module PartialProd(
  input  [15:0] io_multiplicand,
  input  [15:0] io_multiplier,
  output [15:0] io_outs_0,
  output [15:0] io_outs_1,
  output [15:0] io_outs_2,
  output [15:0] io_outs_3,
  output [15:0] io_outs_4,
  output [15:0] io_outs_5,
  output [15:0] io_outs_6,
  output [15:0] io_outs_7,
  output [15:0] io_outs_8,
  output [15:0] io_outs_9,
  output [15:0] io_outs_10,
  output [15:0] io_outs_11,
  output [15:0] io_outs_12,
  output [15:0] io_outs_13,
  output [15:0] io_outs_14,
  output [15:0] io_outs_15
);
  wire  _T_18 = io_multiplicand[0] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_21 = io_multiplicand[1] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_24 = io_multiplicand[2] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_27 = io_multiplicand[3] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_30 = io_multiplicand[4] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_33 = io_multiplicand[5] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_36 = io_multiplicand[6] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_39 = io_multiplicand[7] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_42 = io_multiplicand[8] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_45 = io_multiplicand[9] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_48 = io_multiplicand[10] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_51 = io_multiplicand[11] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_54 = io_multiplicand[12] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_57 = io_multiplicand[13] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_60 = io_multiplicand[14] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_63 = io_multiplicand[15] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire [9:0] _T_72 = {_T_63,_T_60,_T_57,_T_54,_T_51,_T_48,_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58]
  wire [14:0] _T_77 = {_T_72,_T_33,_T_30,_T_27,_T_24,_T_21}; // @[Cat.scala 29:58]
  wire  _T_97 = io_multiplicand[0] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_100 = io_multiplicand[1] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_103 = io_multiplicand[2] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_106 = io_multiplicand[3] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_109 = io_multiplicand[4] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_112 = io_multiplicand[5] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_115 = io_multiplicand[6] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_118 = io_multiplicand[7] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_121 = io_multiplicand[8] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_124 = io_multiplicand[9] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_127 = io_multiplicand[10] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_130 = io_multiplicand[11] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_133 = io_multiplicand[12] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_136 = io_multiplicand[13] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_139 = io_multiplicand[14] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_142 = io_multiplicand[15] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire [9:0] _T_151 = {_T_142,_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118,_T_115}; // @[Cat.scala 29:58]
  wire [14:0] _T_156 = {_T_151,_T_112,_T_109,_T_106,_T_103,_T_100}; // @[Cat.scala 29:58]
  wire  _T_176 = io_multiplicand[0] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_179 = io_multiplicand[1] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_182 = io_multiplicand[2] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_185 = io_multiplicand[3] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_188 = io_multiplicand[4] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_191 = io_multiplicand[5] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_194 = io_multiplicand[6] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_197 = io_multiplicand[7] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_200 = io_multiplicand[8] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_203 = io_multiplicand[9] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_206 = io_multiplicand[10] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_209 = io_multiplicand[11] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_212 = io_multiplicand[12] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_215 = io_multiplicand[13] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_218 = io_multiplicand[14] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_221 = io_multiplicand[15] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire [9:0] _T_230 = {_T_221,_T_218,_T_215,_T_212,_T_209,_T_206,_T_203,_T_200,_T_197,_T_194}; // @[Cat.scala 29:58]
  wire [14:0] _T_235 = {_T_230,_T_191,_T_188,_T_185,_T_182,_T_179}; // @[Cat.scala 29:58]
  wire  _T_255 = io_multiplicand[0] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_258 = io_multiplicand[1] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_261 = io_multiplicand[2] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_264 = io_multiplicand[3] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_267 = io_multiplicand[4] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_270 = io_multiplicand[5] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_273 = io_multiplicand[6] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_276 = io_multiplicand[7] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_279 = io_multiplicand[8] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_282 = io_multiplicand[9] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_285 = io_multiplicand[10] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_288 = io_multiplicand[11] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_291 = io_multiplicand[12] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_294 = io_multiplicand[13] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_297 = io_multiplicand[14] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_300 = io_multiplicand[15] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire [9:0] _T_309 = {_T_300,_T_297,_T_294,_T_291,_T_288,_T_285,_T_282,_T_279,_T_276,_T_273}; // @[Cat.scala 29:58]
  wire [14:0] _T_314 = {_T_309,_T_270,_T_267,_T_264,_T_261,_T_258}; // @[Cat.scala 29:58]
  wire  _T_334 = io_multiplicand[0] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_337 = io_multiplicand[1] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_340 = io_multiplicand[2] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_343 = io_multiplicand[3] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_346 = io_multiplicand[4] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_349 = io_multiplicand[5] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_352 = io_multiplicand[6] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_355 = io_multiplicand[7] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_358 = io_multiplicand[8] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_361 = io_multiplicand[9] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_364 = io_multiplicand[10] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_367 = io_multiplicand[11] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_370 = io_multiplicand[12] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_373 = io_multiplicand[13] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_376 = io_multiplicand[14] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_379 = io_multiplicand[15] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire [9:0] _T_388 = {_T_379,_T_376,_T_373,_T_370,_T_367,_T_364,_T_361,_T_358,_T_355,_T_352}; // @[Cat.scala 29:58]
  wire [14:0] _T_393 = {_T_388,_T_349,_T_346,_T_343,_T_340,_T_337}; // @[Cat.scala 29:58]
  wire  _T_413 = io_multiplicand[0] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_416 = io_multiplicand[1] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_419 = io_multiplicand[2] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_422 = io_multiplicand[3] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_425 = io_multiplicand[4] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_428 = io_multiplicand[5] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_431 = io_multiplicand[6] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_434 = io_multiplicand[7] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_437 = io_multiplicand[8] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_440 = io_multiplicand[9] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_443 = io_multiplicand[10] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_446 = io_multiplicand[11] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_449 = io_multiplicand[12] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_452 = io_multiplicand[13] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_455 = io_multiplicand[14] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_458 = io_multiplicand[15] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire [9:0] _T_467 = {_T_458,_T_455,_T_452,_T_449,_T_446,_T_443,_T_440,_T_437,_T_434,_T_431}; // @[Cat.scala 29:58]
  wire [14:0] _T_472 = {_T_467,_T_428,_T_425,_T_422,_T_419,_T_416}; // @[Cat.scala 29:58]
  wire  _T_492 = io_multiplicand[0] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_495 = io_multiplicand[1] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_498 = io_multiplicand[2] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_501 = io_multiplicand[3] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_504 = io_multiplicand[4] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_507 = io_multiplicand[5] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_510 = io_multiplicand[6] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_513 = io_multiplicand[7] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_516 = io_multiplicand[8] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_519 = io_multiplicand[9] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_522 = io_multiplicand[10] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_525 = io_multiplicand[11] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_528 = io_multiplicand[12] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_531 = io_multiplicand[13] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_534 = io_multiplicand[14] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_537 = io_multiplicand[15] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire [9:0] _T_546 = {_T_537,_T_534,_T_531,_T_528,_T_525,_T_522,_T_519,_T_516,_T_513,_T_510}; // @[Cat.scala 29:58]
  wire [14:0] _T_551 = {_T_546,_T_507,_T_504,_T_501,_T_498,_T_495}; // @[Cat.scala 29:58]
  wire  _T_571 = io_multiplicand[0] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_574 = io_multiplicand[1] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_577 = io_multiplicand[2] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_580 = io_multiplicand[3] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_583 = io_multiplicand[4] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_586 = io_multiplicand[5] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_589 = io_multiplicand[6] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_592 = io_multiplicand[7] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_595 = io_multiplicand[8] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_598 = io_multiplicand[9] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_601 = io_multiplicand[10] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_604 = io_multiplicand[11] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_607 = io_multiplicand[12] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_610 = io_multiplicand[13] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_613 = io_multiplicand[14] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_616 = io_multiplicand[15] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire [9:0] _T_625 = {_T_616,_T_613,_T_610,_T_607,_T_604,_T_601,_T_598,_T_595,_T_592,_T_589}; // @[Cat.scala 29:58]
  wire [14:0] _T_630 = {_T_625,_T_586,_T_583,_T_580,_T_577,_T_574}; // @[Cat.scala 29:58]
  wire  _T_650 = io_multiplicand[0] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_653 = io_multiplicand[1] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_656 = io_multiplicand[2] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_659 = io_multiplicand[3] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_662 = io_multiplicand[4] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_665 = io_multiplicand[5] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_668 = io_multiplicand[6] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_671 = io_multiplicand[7] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_674 = io_multiplicand[8] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_677 = io_multiplicand[9] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_680 = io_multiplicand[10] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_683 = io_multiplicand[11] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_686 = io_multiplicand[12] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_689 = io_multiplicand[13] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_692 = io_multiplicand[14] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_695 = io_multiplicand[15] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire [9:0] _T_704 = {_T_695,_T_692,_T_689,_T_686,_T_683,_T_680,_T_677,_T_674,_T_671,_T_668}; // @[Cat.scala 29:58]
  wire [14:0] _T_709 = {_T_704,_T_665,_T_662,_T_659,_T_656,_T_653}; // @[Cat.scala 29:58]
  wire  _T_729 = io_multiplicand[0] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_732 = io_multiplicand[1] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_735 = io_multiplicand[2] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_738 = io_multiplicand[3] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_741 = io_multiplicand[4] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_744 = io_multiplicand[5] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_747 = io_multiplicand[6] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_750 = io_multiplicand[7] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_753 = io_multiplicand[8] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_756 = io_multiplicand[9] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_759 = io_multiplicand[10] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_762 = io_multiplicand[11] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_765 = io_multiplicand[12] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_768 = io_multiplicand[13] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_771 = io_multiplicand[14] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_774 = io_multiplicand[15] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire [9:0] _T_783 = {_T_774,_T_771,_T_768,_T_765,_T_762,_T_759,_T_756,_T_753,_T_750,_T_747}; // @[Cat.scala 29:58]
  wire [14:0] _T_788 = {_T_783,_T_744,_T_741,_T_738,_T_735,_T_732}; // @[Cat.scala 29:58]
  wire  _T_808 = io_multiplicand[0] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_811 = io_multiplicand[1] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_814 = io_multiplicand[2] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_817 = io_multiplicand[3] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_820 = io_multiplicand[4] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_823 = io_multiplicand[5] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_826 = io_multiplicand[6] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_829 = io_multiplicand[7] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_832 = io_multiplicand[8] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_835 = io_multiplicand[9] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_838 = io_multiplicand[10] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_841 = io_multiplicand[11] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_844 = io_multiplicand[12] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_847 = io_multiplicand[13] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_850 = io_multiplicand[14] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_853 = io_multiplicand[15] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire [9:0] _T_862 = {_T_853,_T_850,_T_847,_T_844,_T_841,_T_838,_T_835,_T_832,_T_829,_T_826}; // @[Cat.scala 29:58]
  wire [14:0] _T_867 = {_T_862,_T_823,_T_820,_T_817,_T_814,_T_811}; // @[Cat.scala 29:58]
  wire  _T_887 = io_multiplicand[0] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_890 = io_multiplicand[1] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_893 = io_multiplicand[2] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_896 = io_multiplicand[3] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_899 = io_multiplicand[4] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_902 = io_multiplicand[5] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_905 = io_multiplicand[6] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_908 = io_multiplicand[7] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_911 = io_multiplicand[8] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_914 = io_multiplicand[9] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_917 = io_multiplicand[10] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_920 = io_multiplicand[11] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_923 = io_multiplicand[12] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_926 = io_multiplicand[13] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_929 = io_multiplicand[14] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_932 = io_multiplicand[15] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire [9:0] _T_941 = {_T_932,_T_929,_T_926,_T_923,_T_920,_T_917,_T_914,_T_911,_T_908,_T_905}; // @[Cat.scala 29:58]
  wire [14:0] _T_946 = {_T_941,_T_902,_T_899,_T_896,_T_893,_T_890}; // @[Cat.scala 29:58]
  wire  _T_966 = io_multiplicand[0] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_969 = io_multiplicand[1] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_972 = io_multiplicand[2] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_975 = io_multiplicand[3] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_978 = io_multiplicand[4] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_981 = io_multiplicand[5] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_984 = io_multiplicand[6] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_987 = io_multiplicand[7] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_990 = io_multiplicand[8] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_993 = io_multiplicand[9] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_996 = io_multiplicand[10] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_999 = io_multiplicand[11] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1002 = io_multiplicand[12] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1005 = io_multiplicand[13] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1008 = io_multiplicand[14] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1011 = io_multiplicand[15] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1020 = {_T_1011,_T_1008,_T_1005,_T_1002,_T_999,_T_996,_T_993,_T_990,_T_987,_T_984}; // @[Cat.scala 29:58]
  wire [14:0] _T_1025 = {_T_1020,_T_981,_T_978,_T_975,_T_972,_T_969}; // @[Cat.scala 29:58]
  wire  _T_1045 = io_multiplicand[0] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1048 = io_multiplicand[1] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1051 = io_multiplicand[2] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1054 = io_multiplicand[3] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1057 = io_multiplicand[4] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1060 = io_multiplicand[5] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1063 = io_multiplicand[6] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1066 = io_multiplicand[7] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1069 = io_multiplicand[8] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1072 = io_multiplicand[9] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1075 = io_multiplicand[10] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1078 = io_multiplicand[11] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1081 = io_multiplicand[12] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1084 = io_multiplicand[13] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1087 = io_multiplicand[14] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1090 = io_multiplicand[15] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1099 = {_T_1090,_T_1087,_T_1084,_T_1081,_T_1078,_T_1075,_T_1072,_T_1069,_T_1066,_T_1063}; // @[Cat.scala 29:58]
  wire [14:0] _T_1104 = {_T_1099,_T_1060,_T_1057,_T_1054,_T_1051,_T_1048}; // @[Cat.scala 29:58]
  wire  _T_1124 = io_multiplicand[0] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1127 = io_multiplicand[1] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1130 = io_multiplicand[2] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1133 = io_multiplicand[3] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1136 = io_multiplicand[4] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1139 = io_multiplicand[5] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1142 = io_multiplicand[6] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1145 = io_multiplicand[7] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1148 = io_multiplicand[8] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1151 = io_multiplicand[9] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1154 = io_multiplicand[10] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1157 = io_multiplicand[11] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1160 = io_multiplicand[12] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1163 = io_multiplicand[13] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1166 = io_multiplicand[14] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1169 = io_multiplicand[15] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1178 = {_T_1169,_T_1166,_T_1163,_T_1160,_T_1157,_T_1154,_T_1151,_T_1148,_T_1145,_T_1142}; // @[Cat.scala 29:58]
  wire [14:0] _T_1183 = {_T_1178,_T_1139,_T_1136,_T_1133,_T_1130,_T_1127}; // @[Cat.scala 29:58]
  wire  _T_1203 = io_multiplicand[0] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1206 = io_multiplicand[1] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1209 = io_multiplicand[2] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1212 = io_multiplicand[3] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1215 = io_multiplicand[4] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1218 = io_multiplicand[5] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1221 = io_multiplicand[6] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1224 = io_multiplicand[7] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1227 = io_multiplicand[8] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1230 = io_multiplicand[9] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1233 = io_multiplicand[10] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1236 = io_multiplicand[11] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1239 = io_multiplicand[12] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1242 = io_multiplicand[13] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1245 = io_multiplicand[14] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1248 = io_multiplicand[15] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1257 = {_T_1248,_T_1245,_T_1242,_T_1239,_T_1236,_T_1233,_T_1230,_T_1227,_T_1224,_T_1221}; // @[Cat.scala 29:58]
  wire [14:0] _T_1262 = {_T_1257,_T_1218,_T_1215,_T_1212,_T_1209,_T_1206}; // @[Cat.scala 29:58]
  assign io_outs_0 = {_T_77,_T_18}; // @[partialprod.scala 18:16]
  assign io_outs_1 = {_T_156,_T_97}; // @[partialprod.scala 18:16]
  assign io_outs_2 = {_T_235,_T_176}; // @[partialprod.scala 18:16]
  assign io_outs_3 = {_T_314,_T_255}; // @[partialprod.scala 18:16]
  assign io_outs_4 = {_T_393,_T_334}; // @[partialprod.scala 18:16]
  assign io_outs_5 = {_T_472,_T_413}; // @[partialprod.scala 18:16]
  assign io_outs_6 = {_T_551,_T_492}; // @[partialprod.scala 18:16]
  assign io_outs_7 = {_T_630,_T_571}; // @[partialprod.scala 18:16]
  assign io_outs_8 = {_T_709,_T_650}; // @[partialprod.scala 18:16]
  assign io_outs_9 = {_T_788,_T_729}; // @[partialprod.scala 18:16]
  assign io_outs_10 = {_T_867,_T_808}; // @[partialprod.scala 18:16]
  assign io_outs_11 = {_T_946,_T_887}; // @[partialprod.scala 18:16]
  assign io_outs_12 = {_T_1025,_T_966}; // @[partialprod.scala 18:16]
  assign io_outs_13 = {_T_1104,_T_1045}; // @[partialprod.scala 18:16]
  assign io_outs_14 = {_T_1183,_T_1124}; // @[partialprod.scala 18:16]
  assign io_outs_15 = {_T_1262,_T_1203}; // @[partialprod.scala 18:16]
endmodule
module FullAdder(
  input   io_a,
  input   io_b,
  input   io_ci,
  output  io_s,
  output  io_co
);
  wire  a_xor_b = io_a ^ io_b; // @[comp.scala 28:22]
  wire  a_and_b = io_a & io_b; // @[comp.scala 31:22]
  wire  a_and_cin = io_a & io_ci; // @[comp.scala 32:24]
  wire  b_and_cin = io_b & io_ci; // @[comp.scala 33:24]
  wire  _T_1 = a_and_b | b_and_cin; // @[comp.scala 34:20]
  assign io_s = a_xor_b ^ io_ci; // @[comp.scala 29:8]
  assign io_co = _T_1 | a_and_cin; // @[comp.scala 34:9]
endmodule
module HalfAdder(
  input   io_a,
  input   io_b,
  output  io_s,
  output  io_co
);
  assign io_s = io_a ^ io_b; // @[comp.scala 15:8]
  assign io_co = io_a & io_b; // @[comp.scala 16:9]
endmodule
module Wallaced(
  input  [15:0] io_pp_0,
  input  [15:0] io_pp_1,
  input  [15:0] io_pp_2,
  input  [15:0] io_pp_3,
  input  [15:0] io_pp_4,
  input  [15:0] io_pp_5,
  input  [15:0] io_pp_6,
  input  [15:0] io_pp_7,
  input  [15:0] io_pp_8,
  input  [15:0] io_pp_9,
  input  [15:0] io_pp_10,
  input  [15:0] io_pp_11,
  input  [15:0] io_pp_12,
  input  [15:0] io_pp_13,
  input  [15:0] io_pp_14,
  input  [15:0] io_pp_15,
  input  [15:0] io_pp_16,
  input  [15:0] io_pp_17,
  input  [15:0] io_pp_18,
  input  [15:0] io_pp_19,
  input  [15:0] io_pp_20,
  input  [15:0] io_pp_21,
  input  [15:0] io_pp_22,
  input  [15:0] io_pp_23,
  input  [15:0] io_pp_24,
  input  [15:0] io_pp_25,
  input  [15:0] io_pp_26,
  input  [15:0] io_pp_27,
  input  [15:0] io_pp_28,
  input  [15:0] io_pp_29,
  input  [15:0] io_pp_30,
  input  [15:0] io_pp_31,
  output [31:0] io_augend,
  output [31:0] io_addend
);
  wire  FullAdder_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_1_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_1_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_1_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_1_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_1_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_2_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_2_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_2_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_2_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_2_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_3_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_3_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_3_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_3_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_3_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_4_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_4_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_4_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_4_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_4_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_5_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_5_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_5_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_5_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_5_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_6_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_6_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_6_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_6_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_6_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_7_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_7_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_7_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_7_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_7_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_8_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_8_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_8_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_8_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_8_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_9_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_9_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_9_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_9_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_9_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_10_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_10_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_10_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_10_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_10_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_11_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_11_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_11_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_11_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_11_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_12_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_12_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_12_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_12_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_12_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_13_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_13_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_13_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_13_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_13_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_14_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_14_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_14_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_14_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_14_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_15_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_15_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_15_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_15_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_15_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_16_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_16_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_16_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_16_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_16_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_17_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_17_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_17_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_17_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_17_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_18_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_18_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_18_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_18_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_18_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_19_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_19_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_19_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_19_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_19_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_20_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_20_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_20_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_20_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_20_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_21_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_21_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_21_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_21_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_21_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_22_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_22_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_22_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_22_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_22_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_23_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_23_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_23_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_23_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_23_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_24_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_24_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_24_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_24_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_24_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_25_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_25_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_25_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_25_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_25_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_26_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_26_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_26_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_26_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_26_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_27_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_27_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_27_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_27_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_27_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_28_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_28_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_28_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_28_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_28_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_29_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_29_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_29_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_29_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_29_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_30_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_30_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_30_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_30_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_30_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_31_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_31_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_31_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_31_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_31_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_32_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_32_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_32_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_32_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_32_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_33_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_33_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_33_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_33_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_33_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_34_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_34_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_34_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_34_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_34_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_35_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_35_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_35_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_35_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_35_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_36_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_36_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_36_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_36_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_36_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_37_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_37_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_37_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_37_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_37_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_38_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_38_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_38_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_38_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_38_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_39_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_39_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_39_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_39_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_39_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_40_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_40_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_40_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_40_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_40_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_41_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_41_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_41_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_41_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_41_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_42_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_42_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_42_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_42_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_42_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_43_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_43_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_43_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_43_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_43_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_44_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_44_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_44_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_44_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_44_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_45_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_45_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_45_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_45_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_45_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_46_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_46_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_46_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_46_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_46_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_47_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_47_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_47_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_47_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_47_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_48_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_48_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_48_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_48_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_48_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_49_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_49_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_49_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_49_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_49_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_50_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_50_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_50_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_50_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_50_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_51_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_51_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_51_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_51_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_51_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_52_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_52_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_52_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_52_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_52_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_53_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_53_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_53_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_53_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_53_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_54_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_54_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_54_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_54_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_54_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_55_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_55_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_55_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_55_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_55_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_56_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_56_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_56_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_56_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_56_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_57_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_57_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_57_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_57_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_57_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_58_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_58_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_58_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_58_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_58_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_59_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_59_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_59_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_59_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_59_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_60_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_60_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_60_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_60_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_60_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_61_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_61_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_61_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_61_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_61_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_62_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_62_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_62_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_62_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_62_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_63_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_63_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_63_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_63_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_63_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_64_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_64_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_64_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_64_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_64_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_65_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_65_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_65_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_65_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_65_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_66_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_66_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_66_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_66_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_66_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_67_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_67_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_67_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_67_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_67_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_68_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_68_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_68_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_68_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_68_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_69_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_69_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_69_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_69_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_69_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_70_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_70_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_70_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_70_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_70_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_71_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_71_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_71_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_71_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_71_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_72_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_72_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_72_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_72_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_72_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_73_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_73_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_73_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_73_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_73_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_74_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_74_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_74_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_74_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_74_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_75_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_75_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_75_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_75_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_75_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_76_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_76_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_76_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_76_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_76_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_77_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_77_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_77_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_77_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_77_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_78_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_78_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_78_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_78_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_78_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_79_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_79_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_79_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_79_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_79_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_80_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_80_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_80_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_80_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_80_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_81_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_81_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_81_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_81_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_81_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_82_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_82_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_82_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_82_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_82_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_83_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_83_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_83_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_83_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_83_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_84_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_84_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_84_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_84_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_84_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_85_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_85_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_85_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_85_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_85_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_86_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_86_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_86_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_86_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_86_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_87_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_87_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_87_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_87_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_87_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_88_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_88_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_88_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_88_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_88_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_89_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_89_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_89_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_89_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_89_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_90_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_90_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_90_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_90_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_90_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_91_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_91_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_91_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_91_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_91_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_92_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_92_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_92_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_92_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_92_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_93_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_93_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_93_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_93_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_93_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_94_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_94_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_94_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_94_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_94_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_95_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_95_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_95_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_95_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_95_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_96_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_96_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_96_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_96_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_96_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_97_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_97_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_97_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_97_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_97_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_98_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_98_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_98_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_98_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_98_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_99_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_99_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_99_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_99_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_99_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_100_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_100_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_100_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_100_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_100_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_101_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_101_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_101_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_101_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_101_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_102_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_102_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_102_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_102_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_102_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_103_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_103_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_103_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_103_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_103_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_104_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_104_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_104_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_104_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_104_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_105_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_105_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_105_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_105_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_105_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_106_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_106_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_106_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_106_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_106_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_107_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_107_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_107_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_107_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_107_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_108_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_108_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_108_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_108_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_108_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_109_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_109_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_109_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_109_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_109_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_110_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_110_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_110_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_110_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_110_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_111_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_111_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_111_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_111_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_111_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_112_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_112_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_112_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_112_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_112_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_113_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_113_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_113_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_113_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_113_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_114_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_114_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_114_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_114_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_114_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_115_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_115_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_115_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_115_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_115_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_116_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_116_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_116_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_116_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_116_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_117_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_117_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_117_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_117_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_117_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_118_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_118_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_118_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_118_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_118_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_119_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_119_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_119_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_119_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_119_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_120_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_120_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_120_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_120_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_120_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_121_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_121_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_121_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_121_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_121_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_122_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_122_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_122_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_122_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_122_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_123_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_123_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_123_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_123_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_123_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_124_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_124_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_124_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_124_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_124_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_125_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_125_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_125_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_125_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_125_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_126_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_126_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_126_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_126_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_126_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_127_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_127_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_127_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_127_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_127_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_128_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_128_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_128_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_128_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_128_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_129_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_129_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_129_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_129_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_129_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_130_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_130_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_130_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_130_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_130_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_131_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_131_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_131_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_131_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_131_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_132_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_132_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_132_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_132_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_132_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_133_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_133_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_133_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_133_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_133_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_134_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_134_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_134_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_134_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_134_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_135_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_135_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_135_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_135_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_135_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_136_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_136_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_136_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_136_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_136_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_137_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_137_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_137_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_137_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_137_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_138_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_138_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_138_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_138_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_138_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_139_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_139_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_139_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_139_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_139_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_140_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_140_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_140_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_140_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_140_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_141_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_141_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_141_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_141_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_141_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_142_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_142_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_142_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_142_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_142_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_143_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_143_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_143_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_143_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_143_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_144_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_144_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_144_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_144_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_144_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_145_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_145_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_145_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_145_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_145_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_146_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_146_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_146_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_146_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_146_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_147_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_147_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_147_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_147_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_147_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_148_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_148_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_148_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_148_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_148_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_149_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_149_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_149_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_149_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_149_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_150_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_150_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_150_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_150_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_150_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_151_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_151_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_151_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_151_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_151_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_152_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_152_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_152_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_152_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_152_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_153_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_153_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_153_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_153_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_153_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_154_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_154_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_154_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_154_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_154_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_155_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_155_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_155_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_155_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_155_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_156_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_156_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_156_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_156_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_156_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_157_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_157_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_157_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_157_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_157_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_158_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_158_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_158_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_158_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_158_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_159_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_159_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_159_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_159_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_159_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_160_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_160_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_160_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_160_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_160_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_161_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_161_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_161_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_161_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_161_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_162_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_162_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_162_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_162_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_162_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_163_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_163_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_163_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_163_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_163_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_164_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_164_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_164_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_164_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_164_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_165_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_165_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_165_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_165_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_165_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_166_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_166_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_166_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_166_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_166_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_167_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_167_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_167_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_167_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_167_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_168_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_168_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_168_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_168_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_168_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_169_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_169_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_169_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_169_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_169_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_170_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_170_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_170_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_170_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_170_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_171_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_171_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_171_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_171_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_171_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_172_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_172_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_172_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_172_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_172_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_173_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_173_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_173_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_173_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_173_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_174_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_174_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_174_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_174_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_174_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_1_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_1_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_1_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_1_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_175_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_175_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_175_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_175_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_175_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_176_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_176_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_176_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_176_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_176_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_177_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_177_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_177_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_177_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_177_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_178_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_178_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_178_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_178_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_178_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_179_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_179_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_179_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_179_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_179_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_180_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_180_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_180_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_180_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_180_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_181_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_181_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_181_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_181_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_181_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_182_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_182_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_182_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_182_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_182_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_183_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_183_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_183_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_183_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_183_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_184_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_184_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_184_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_184_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_184_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_185_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_185_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_185_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_185_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_185_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_186_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_186_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_186_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_186_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_186_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_187_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_187_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_187_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_187_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_187_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_2_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_2_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_2_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_2_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_188_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_188_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_188_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_188_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_188_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_189_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_189_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_189_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_189_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_189_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_190_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_190_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_190_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_190_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_190_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_191_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_191_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_191_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_191_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_191_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_192_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_192_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_192_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_192_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_192_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_193_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_193_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_193_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_193_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_193_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_194_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_194_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_194_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_194_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_194_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_195_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_195_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_195_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_195_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_195_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_196_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_196_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_196_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_196_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_196_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_197_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_197_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_197_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_197_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_197_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_198_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_198_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_198_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_198_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_198_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_199_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_199_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_199_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_199_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_199_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_200_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_200_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_200_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_200_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_200_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_3_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_3_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_3_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_3_io_co; // @[wallaced.scala 77:25]
  wire  HalfAdder_4_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_4_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_4_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_4_io_co; // @[wallaced.scala 77:25]
  wire  HalfAdder_5_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_5_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_5_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_5_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_201_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_201_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_201_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_201_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_201_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_202_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_202_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_202_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_202_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_202_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_203_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_203_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_203_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_203_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_203_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_204_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_204_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_204_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_204_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_204_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_205_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_205_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_205_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_205_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_205_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_206_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_206_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_206_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_206_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_206_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_207_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_207_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_207_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_207_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_207_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_208_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_208_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_208_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_208_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_208_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_209_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_209_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_209_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_209_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_209_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_210_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_210_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_210_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_210_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_210_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_211_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_211_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_211_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_211_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_211_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_212_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_212_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_212_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_212_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_212_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_213_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_213_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_213_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_213_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_213_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_214_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_214_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_214_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_214_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_214_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_215_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_215_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_215_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_215_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_215_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_216_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_216_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_216_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_216_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_216_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_217_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_217_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_217_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_217_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_217_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_218_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_218_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_218_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_218_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_218_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_219_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_219_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_219_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_219_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_219_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_220_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_220_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_220_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_220_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_220_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_221_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_221_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_221_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_221_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_221_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_222_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_222_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_222_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_222_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_222_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_223_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_223_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_223_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_223_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_223_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_224_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_224_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_224_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_224_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_224_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_225_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_225_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_225_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_225_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_225_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_226_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_226_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_226_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_226_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_226_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_227_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_227_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_227_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_227_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_227_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_228_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_228_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_228_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_228_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_228_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_229_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_229_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_229_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_229_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_229_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_230_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_230_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_230_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_230_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_230_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_231_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_231_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_231_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_231_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_231_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_232_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_232_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_232_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_232_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_232_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_233_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_233_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_233_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_233_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_233_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_234_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_234_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_234_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_234_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_234_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_235_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_235_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_235_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_235_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_235_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_236_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_236_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_236_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_236_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_236_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_237_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_237_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_237_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_237_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_237_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_238_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_238_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_238_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_238_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_238_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_239_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_239_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_239_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_239_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_239_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_240_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_240_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_240_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_240_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_240_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_241_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_241_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_241_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_241_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_241_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_242_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_242_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_242_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_242_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_242_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_243_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_243_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_243_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_243_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_243_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_244_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_244_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_244_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_244_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_244_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_245_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_245_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_245_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_245_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_245_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_246_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_246_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_246_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_246_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_246_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_247_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_247_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_247_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_247_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_247_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_248_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_248_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_248_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_248_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_248_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_249_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_249_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_249_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_249_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_249_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_250_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_250_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_250_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_250_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_250_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_251_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_251_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_251_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_251_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_251_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_252_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_252_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_252_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_252_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_252_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_253_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_253_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_253_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_253_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_253_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_254_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_254_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_254_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_254_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_254_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_255_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_255_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_255_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_255_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_255_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_256_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_256_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_256_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_256_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_256_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_257_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_257_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_257_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_257_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_257_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_258_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_258_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_258_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_258_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_258_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_259_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_259_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_259_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_259_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_259_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_260_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_260_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_260_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_260_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_260_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_261_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_261_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_261_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_261_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_261_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_262_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_262_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_262_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_262_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_262_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_263_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_263_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_263_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_263_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_263_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_264_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_264_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_264_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_264_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_264_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_265_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_265_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_265_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_265_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_265_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_266_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_266_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_266_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_266_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_266_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_267_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_267_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_267_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_267_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_267_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_268_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_268_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_268_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_268_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_268_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_269_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_269_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_269_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_269_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_269_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_270_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_270_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_270_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_270_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_270_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_271_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_271_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_271_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_271_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_271_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_272_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_272_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_272_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_272_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_272_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_273_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_273_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_273_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_273_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_273_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_274_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_274_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_274_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_274_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_274_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_275_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_275_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_275_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_275_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_275_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_276_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_276_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_276_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_276_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_276_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_277_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_277_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_277_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_277_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_277_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_278_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_278_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_278_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_278_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_278_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_279_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_279_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_279_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_279_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_279_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_280_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_280_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_280_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_280_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_280_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_281_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_281_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_281_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_281_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_281_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_282_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_282_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_282_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_282_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_282_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_283_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_283_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_283_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_283_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_283_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_284_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_284_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_284_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_284_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_284_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_285_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_285_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_285_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_285_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_285_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_286_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_286_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_286_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_286_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_286_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_287_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_287_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_287_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_287_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_287_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_288_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_288_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_288_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_288_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_288_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_289_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_289_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_289_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_289_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_289_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_290_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_290_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_290_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_290_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_290_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_291_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_291_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_291_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_291_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_291_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_292_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_292_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_292_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_292_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_292_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_293_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_293_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_293_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_293_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_293_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_294_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_294_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_294_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_294_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_294_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_295_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_295_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_295_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_295_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_295_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_296_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_296_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_296_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_296_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_296_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_297_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_297_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_297_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_297_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_297_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_298_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_298_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_298_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_298_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_298_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_299_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_299_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_299_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_299_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_299_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_300_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_300_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_300_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_300_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_300_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_301_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_301_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_301_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_301_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_301_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_302_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_302_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_302_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_302_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_302_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_303_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_303_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_303_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_303_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_303_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_304_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_304_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_304_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_304_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_304_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_305_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_305_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_305_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_305_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_305_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_306_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_306_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_306_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_306_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_306_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_307_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_307_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_307_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_307_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_307_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_308_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_308_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_308_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_308_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_308_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_309_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_309_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_309_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_309_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_309_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_310_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_310_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_310_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_310_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_310_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_311_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_311_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_311_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_311_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_311_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_312_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_312_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_312_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_312_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_312_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_313_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_313_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_313_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_313_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_313_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_314_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_314_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_314_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_314_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_314_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_315_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_315_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_315_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_315_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_315_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_316_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_316_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_316_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_316_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_316_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_317_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_317_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_317_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_317_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_317_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_318_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_318_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_318_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_318_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_318_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_319_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_319_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_319_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_319_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_319_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_320_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_320_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_320_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_320_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_320_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_321_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_321_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_321_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_321_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_321_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_322_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_322_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_322_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_322_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_322_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_323_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_323_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_323_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_323_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_323_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_324_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_324_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_324_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_324_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_324_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_325_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_325_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_325_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_325_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_325_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_326_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_326_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_326_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_326_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_326_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_327_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_327_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_327_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_327_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_327_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_328_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_328_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_328_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_328_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_328_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_329_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_329_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_329_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_329_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_329_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_330_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_330_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_330_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_330_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_330_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_331_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_331_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_331_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_331_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_331_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_332_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_332_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_332_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_332_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_332_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_333_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_333_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_333_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_333_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_333_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_334_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_334_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_334_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_334_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_334_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_335_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_335_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_335_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_335_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_335_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_336_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_336_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_336_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_336_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_336_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_337_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_337_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_337_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_337_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_337_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_338_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_338_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_338_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_338_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_338_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_339_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_339_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_339_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_339_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_339_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_340_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_340_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_340_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_340_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_340_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_341_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_341_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_341_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_341_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_341_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_342_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_342_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_342_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_342_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_342_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_343_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_343_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_343_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_343_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_343_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_344_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_344_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_344_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_344_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_344_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_345_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_345_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_345_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_345_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_345_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_346_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_346_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_346_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_346_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_346_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_347_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_347_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_347_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_347_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_347_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_348_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_348_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_348_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_348_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_348_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_349_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_349_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_349_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_349_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_349_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_350_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_350_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_350_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_350_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_350_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_351_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_351_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_351_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_351_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_351_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_352_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_352_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_352_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_352_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_352_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_353_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_353_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_353_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_353_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_353_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_354_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_354_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_354_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_354_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_354_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_355_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_355_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_355_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_355_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_355_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_356_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_356_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_356_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_356_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_356_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_357_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_357_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_357_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_357_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_357_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_6_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_6_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_6_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_6_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_358_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_358_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_358_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_358_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_358_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_359_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_359_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_359_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_359_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_359_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_360_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_360_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_360_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_360_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_360_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_361_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_361_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_361_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_361_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_361_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_362_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_362_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_362_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_362_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_362_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_363_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_363_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_363_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_363_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_363_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_364_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_364_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_364_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_364_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_364_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_365_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_365_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_365_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_365_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_365_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_366_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_366_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_366_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_366_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_366_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_367_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_367_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_367_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_367_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_367_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_368_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_368_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_368_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_368_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_368_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_369_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_369_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_369_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_369_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_369_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_370_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_370_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_370_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_370_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_370_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_371_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_371_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_371_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_371_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_371_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_372_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_372_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_372_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_372_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_372_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_373_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_373_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_373_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_373_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_373_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_374_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_374_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_374_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_374_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_374_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_375_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_375_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_375_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_375_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_375_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_376_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_376_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_376_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_376_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_376_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_377_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_377_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_377_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_377_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_377_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_378_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_378_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_378_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_378_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_378_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_7_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_7_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_7_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_7_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_379_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_379_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_379_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_379_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_379_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_380_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_380_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_380_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_380_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_380_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_381_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_381_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_381_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_381_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_381_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_382_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_382_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_382_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_382_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_382_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_383_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_383_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_383_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_383_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_383_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_384_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_384_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_384_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_384_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_384_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_385_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_385_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_385_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_385_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_385_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_386_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_386_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_386_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_386_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_386_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_387_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_387_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_387_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_387_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_387_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_388_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_388_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_388_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_388_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_388_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_389_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_389_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_389_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_389_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_389_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_390_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_390_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_390_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_390_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_390_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_391_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_391_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_391_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_391_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_391_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_8_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_8_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_8_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_8_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_392_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_392_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_392_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_392_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_392_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_393_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_393_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_393_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_393_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_393_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_394_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_394_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_394_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_394_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_394_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_395_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_395_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_395_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_395_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_395_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_396_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_396_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_396_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_396_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_396_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_397_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_397_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_397_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_397_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_397_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_398_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_398_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_398_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_398_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_398_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_399_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_399_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_399_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_399_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_399_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_400_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_400_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_400_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_400_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_400_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_401_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_401_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_401_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_401_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_401_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_402_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_402_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_402_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_402_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_402_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_403_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_403_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_403_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_403_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_403_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_404_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_404_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_404_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_404_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_404_io_co; // @[wallaced.scala 86:25]
  wire  HalfAdder_9_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_9_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_9_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_9_io_co; // @[wallaced.scala 77:25]
  wire  HalfAdder_10_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_10_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_10_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_10_io_co; // @[wallaced.scala 77:25]
  wire  HalfAdder_11_io_a; // @[wallaced.scala 77:25]
  wire  HalfAdder_11_io_b; // @[wallaced.scala 77:25]
  wire  HalfAdder_11_io_s; // @[wallaced.scala 77:25]
  wire  HalfAdder_11_io_co; // @[wallaced.scala 77:25]
  wire  FullAdder_405_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_405_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_405_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_405_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_405_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_406_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_406_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_406_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_406_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_406_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_407_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_407_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_407_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_407_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_407_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_408_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_408_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_408_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_408_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_408_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_409_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_409_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_409_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_409_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_409_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_410_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_410_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_410_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_410_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_410_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_411_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_411_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_411_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_411_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_411_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_412_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_412_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_412_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_412_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_412_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_413_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_413_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_413_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_413_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_413_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_414_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_414_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_414_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_414_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_414_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_415_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_415_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_415_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_415_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_415_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_416_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_416_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_416_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_416_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_416_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_417_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_417_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_417_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_417_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_417_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_418_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_418_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_418_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_418_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_418_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_419_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_419_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_419_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_419_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_419_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_420_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_420_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_420_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_420_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_420_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_421_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_421_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_421_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_421_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_421_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_422_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_422_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_422_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_422_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_422_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_423_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_423_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_423_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_423_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_423_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_424_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_424_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_424_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_424_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_424_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_425_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_425_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_425_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_425_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_425_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_426_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_426_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_426_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_426_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_426_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_427_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_427_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_427_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_427_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_427_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_428_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_428_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_428_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_428_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_428_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_429_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_429_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_429_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_429_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_429_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_430_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_430_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_430_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_430_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_430_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_431_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_431_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_431_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_431_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_431_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_432_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_432_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_432_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_432_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_432_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_433_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_433_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_433_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_433_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_433_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_434_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_434_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_434_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_434_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_434_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_435_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_435_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_435_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_435_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_435_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_436_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_436_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_436_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_436_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_436_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_437_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_437_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_437_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_437_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_437_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_438_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_438_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_438_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_438_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_438_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_439_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_439_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_439_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_439_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_439_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_440_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_440_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_440_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_440_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_440_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_441_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_441_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_441_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_441_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_441_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_442_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_442_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_442_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_442_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_442_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_443_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_443_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_443_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_443_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_443_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_444_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_444_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_444_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_444_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_444_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_445_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_445_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_445_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_445_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_445_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_446_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_446_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_446_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_446_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_446_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_447_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_447_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_447_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_447_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_447_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_448_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_448_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_448_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_448_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_448_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_449_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_449_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_449_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_449_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_449_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_450_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_450_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_450_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_450_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_450_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_451_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_451_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_451_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_451_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_451_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_452_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_452_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_452_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_452_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_452_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_453_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_453_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_453_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_453_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_453_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_454_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_454_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_454_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_454_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_454_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_455_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_455_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_455_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_455_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_455_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_456_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_456_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_456_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_456_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_456_io_co; // @[wallaced.scala 86:25]
  wire  FullAdder_457_io_a; // @[wallaced.scala 86:25]
  wire  FullAdder_457_io_b; // @[wallaced.scala 86:25]
  wire  FullAdder_457_io_ci; // @[wallaced.scala 86:25]
  wire  FullAdder_457_io_s; // @[wallaced.scala 86:25]
  wire  FullAdder_457_io_co; // @[wallaced.scala 86:25]
  wire  res0_0 = io_pp_0[0]; // @[wallaced.scala 56:49]
  wire  res1_0 = io_pp_16[0]; // @[wallaced.scala 56:49]
  wire  res0_1 = io_pp_17[0]; // @[wallaced.scala 56:49]
  wire  res0_31 = FullAdder_408_io_co; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_30 = FullAdder_429_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_29 = FullAdder_430_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_28 = FullAdder_431_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_27 = FullAdder_432_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_26 = FullAdder_433_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_25 = FullAdder_434_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_24 = FullAdder_435_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_23 = FullAdder_436_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_22 = FullAdder_437_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire [9:0] _T_520 = {res0_31,res0_30,res0_29,res0_28,res0_27,res0_26,res0_25,res0_24,res0_23,res0_22}; // @[Cat.scala 29:58]
  wire  res0_21 = FullAdder_438_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_20 = FullAdder_439_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_19 = FullAdder_440_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_18 = FullAdder_441_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_17 = FullAdder_442_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_16 = FullAdder_443_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_15 = FullAdder_444_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_14 = FullAdder_445_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_13 = FullAdder_449_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire [18:0] _T_529 = {_T_520,res0_21,res0_20,res0_19,res0_18,res0_17,res0_16,res0_15,res0_14,res0_13}; // @[Cat.scala 29:58]
  wire  res0_12 = FullAdder_446_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_11 = FullAdder_453_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_10 = FullAdder_450_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_9 = FullAdder_447_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_8 = FullAdder_457_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_7 = FullAdder_456_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_6 = FullAdder_455_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_5 = FullAdder_454_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_4 = FullAdder_452_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire [27:0] _T_538 = {_T_529,res0_12,res0_11,res0_10,res0_9,res0_8,res0_7,res0_6,res0_5,res0_4}; // @[Cat.scala 29:58]
  wire  res0_3 = FullAdder_451_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire  res0_2 = FullAdder_448_io_s; // @[wallaced.scala 97:49 wallaced.scala 102:13]
  wire [30:0] _T_541 = {_T_538,res0_3,res0_2,res0_1}; // @[Cat.scala 29:58]
  wire  res1_31 = FullAdder_429_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_30 = FullAdder_430_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_29 = FullAdder_431_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_28 = FullAdder_432_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_27 = FullAdder_433_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_26 = FullAdder_434_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_25 = FullAdder_435_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_24 = FullAdder_436_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_23 = FullAdder_437_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_22 = FullAdder_438_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire [9:0] _T_551 = {res1_31,res1_30,res1_29,res1_28,res1_27,res1_26,res1_25,res1_24,res1_23,res1_22}; // @[Cat.scala 29:58]
  wire  res1_21 = FullAdder_439_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_20 = FullAdder_440_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_19 = FullAdder_441_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_18 = FullAdder_442_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_17 = FullAdder_443_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_16 = FullAdder_444_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_15 = FullAdder_445_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_14 = FullAdder_449_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire [18:0] _T_560 = {_T_551,res1_21,res1_20,res1_19,res1_18,res1_17,res1_16,res1_15,res1_14,1'h0}; // @[Cat.scala 29:58]
  wire  res1_12 = FullAdder_453_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire  res1_9 = FullAdder_457_io_co; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire [27:0] _T_569 = {_T_560,res1_12,1'h0,1'h0,res1_9,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire  res1_1 = FullAdder_428_io_s; // @[wallaced.scala 98:49 wallaced.scala 106:15]
  wire [30:0] _T_572 = {_T_569,1'h0,1'h0,res1_1}; // @[Cat.scala 29:58]
  FullAdder FullAdder ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_io_a),
    .io_b(FullAdder_io_b),
    .io_ci(FullAdder_io_ci),
    .io_s(FullAdder_io_s),
    .io_co(FullAdder_io_co)
  );
  FullAdder FullAdder_1 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_1_io_a),
    .io_b(FullAdder_1_io_b),
    .io_ci(FullAdder_1_io_ci),
    .io_s(FullAdder_1_io_s),
    .io_co(FullAdder_1_io_co)
  );
  FullAdder FullAdder_2 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_2_io_a),
    .io_b(FullAdder_2_io_b),
    .io_ci(FullAdder_2_io_ci),
    .io_s(FullAdder_2_io_s),
    .io_co(FullAdder_2_io_co)
  );
  FullAdder FullAdder_3 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_3_io_a),
    .io_b(FullAdder_3_io_b),
    .io_ci(FullAdder_3_io_ci),
    .io_s(FullAdder_3_io_s),
    .io_co(FullAdder_3_io_co)
  );
  FullAdder FullAdder_4 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_4_io_a),
    .io_b(FullAdder_4_io_b),
    .io_ci(FullAdder_4_io_ci),
    .io_s(FullAdder_4_io_s),
    .io_co(FullAdder_4_io_co)
  );
  FullAdder FullAdder_5 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_5_io_a),
    .io_b(FullAdder_5_io_b),
    .io_ci(FullAdder_5_io_ci),
    .io_s(FullAdder_5_io_s),
    .io_co(FullAdder_5_io_co)
  );
  FullAdder FullAdder_6 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_6_io_a),
    .io_b(FullAdder_6_io_b),
    .io_ci(FullAdder_6_io_ci),
    .io_s(FullAdder_6_io_s),
    .io_co(FullAdder_6_io_co)
  );
  FullAdder FullAdder_7 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_7_io_a),
    .io_b(FullAdder_7_io_b),
    .io_ci(FullAdder_7_io_ci),
    .io_s(FullAdder_7_io_s),
    .io_co(FullAdder_7_io_co)
  );
  FullAdder FullAdder_8 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_8_io_a),
    .io_b(FullAdder_8_io_b),
    .io_ci(FullAdder_8_io_ci),
    .io_s(FullAdder_8_io_s),
    .io_co(FullAdder_8_io_co)
  );
  FullAdder FullAdder_9 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_9_io_a),
    .io_b(FullAdder_9_io_b),
    .io_ci(FullAdder_9_io_ci),
    .io_s(FullAdder_9_io_s),
    .io_co(FullAdder_9_io_co)
  );
  FullAdder FullAdder_10 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_10_io_a),
    .io_b(FullAdder_10_io_b),
    .io_ci(FullAdder_10_io_ci),
    .io_s(FullAdder_10_io_s),
    .io_co(FullAdder_10_io_co)
  );
  FullAdder FullAdder_11 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_11_io_a),
    .io_b(FullAdder_11_io_b),
    .io_ci(FullAdder_11_io_ci),
    .io_s(FullAdder_11_io_s),
    .io_co(FullAdder_11_io_co)
  );
  FullAdder FullAdder_12 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_12_io_a),
    .io_b(FullAdder_12_io_b),
    .io_ci(FullAdder_12_io_ci),
    .io_s(FullAdder_12_io_s),
    .io_co(FullAdder_12_io_co)
  );
  FullAdder FullAdder_13 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_13_io_a),
    .io_b(FullAdder_13_io_b),
    .io_ci(FullAdder_13_io_ci),
    .io_s(FullAdder_13_io_s),
    .io_co(FullAdder_13_io_co)
  );
  FullAdder FullAdder_14 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_14_io_a),
    .io_b(FullAdder_14_io_b),
    .io_ci(FullAdder_14_io_ci),
    .io_s(FullAdder_14_io_s),
    .io_co(FullAdder_14_io_co)
  );
  FullAdder FullAdder_15 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_15_io_a),
    .io_b(FullAdder_15_io_b),
    .io_ci(FullAdder_15_io_ci),
    .io_s(FullAdder_15_io_s),
    .io_co(FullAdder_15_io_co)
  );
  FullAdder FullAdder_16 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_16_io_a),
    .io_b(FullAdder_16_io_b),
    .io_ci(FullAdder_16_io_ci),
    .io_s(FullAdder_16_io_s),
    .io_co(FullAdder_16_io_co)
  );
  FullAdder FullAdder_17 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_17_io_a),
    .io_b(FullAdder_17_io_b),
    .io_ci(FullAdder_17_io_ci),
    .io_s(FullAdder_17_io_s),
    .io_co(FullAdder_17_io_co)
  );
  FullAdder FullAdder_18 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_18_io_a),
    .io_b(FullAdder_18_io_b),
    .io_ci(FullAdder_18_io_ci),
    .io_s(FullAdder_18_io_s),
    .io_co(FullAdder_18_io_co)
  );
  FullAdder FullAdder_19 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_19_io_a),
    .io_b(FullAdder_19_io_b),
    .io_ci(FullAdder_19_io_ci),
    .io_s(FullAdder_19_io_s),
    .io_co(FullAdder_19_io_co)
  );
  FullAdder FullAdder_20 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_20_io_a),
    .io_b(FullAdder_20_io_b),
    .io_ci(FullAdder_20_io_ci),
    .io_s(FullAdder_20_io_s),
    .io_co(FullAdder_20_io_co)
  );
  FullAdder FullAdder_21 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_21_io_a),
    .io_b(FullAdder_21_io_b),
    .io_ci(FullAdder_21_io_ci),
    .io_s(FullAdder_21_io_s),
    .io_co(FullAdder_21_io_co)
  );
  FullAdder FullAdder_22 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_22_io_a),
    .io_b(FullAdder_22_io_b),
    .io_ci(FullAdder_22_io_ci),
    .io_s(FullAdder_22_io_s),
    .io_co(FullAdder_22_io_co)
  );
  FullAdder FullAdder_23 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_23_io_a),
    .io_b(FullAdder_23_io_b),
    .io_ci(FullAdder_23_io_ci),
    .io_s(FullAdder_23_io_s),
    .io_co(FullAdder_23_io_co)
  );
  FullAdder FullAdder_24 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_24_io_a),
    .io_b(FullAdder_24_io_b),
    .io_ci(FullAdder_24_io_ci),
    .io_s(FullAdder_24_io_s),
    .io_co(FullAdder_24_io_co)
  );
  FullAdder FullAdder_25 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_25_io_a),
    .io_b(FullAdder_25_io_b),
    .io_ci(FullAdder_25_io_ci),
    .io_s(FullAdder_25_io_s),
    .io_co(FullAdder_25_io_co)
  );
  FullAdder FullAdder_26 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_26_io_a),
    .io_b(FullAdder_26_io_b),
    .io_ci(FullAdder_26_io_ci),
    .io_s(FullAdder_26_io_s),
    .io_co(FullAdder_26_io_co)
  );
  FullAdder FullAdder_27 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_27_io_a),
    .io_b(FullAdder_27_io_b),
    .io_ci(FullAdder_27_io_ci),
    .io_s(FullAdder_27_io_s),
    .io_co(FullAdder_27_io_co)
  );
  FullAdder FullAdder_28 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_28_io_a),
    .io_b(FullAdder_28_io_b),
    .io_ci(FullAdder_28_io_ci),
    .io_s(FullAdder_28_io_s),
    .io_co(FullAdder_28_io_co)
  );
  FullAdder FullAdder_29 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_29_io_a),
    .io_b(FullAdder_29_io_b),
    .io_ci(FullAdder_29_io_ci),
    .io_s(FullAdder_29_io_s),
    .io_co(FullAdder_29_io_co)
  );
  FullAdder FullAdder_30 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_30_io_a),
    .io_b(FullAdder_30_io_b),
    .io_ci(FullAdder_30_io_ci),
    .io_s(FullAdder_30_io_s),
    .io_co(FullAdder_30_io_co)
  );
  FullAdder FullAdder_31 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_31_io_a),
    .io_b(FullAdder_31_io_b),
    .io_ci(FullAdder_31_io_ci),
    .io_s(FullAdder_31_io_s),
    .io_co(FullAdder_31_io_co)
  );
  FullAdder FullAdder_32 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_32_io_a),
    .io_b(FullAdder_32_io_b),
    .io_ci(FullAdder_32_io_ci),
    .io_s(FullAdder_32_io_s),
    .io_co(FullAdder_32_io_co)
  );
  FullAdder FullAdder_33 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_33_io_a),
    .io_b(FullAdder_33_io_b),
    .io_ci(FullAdder_33_io_ci),
    .io_s(FullAdder_33_io_s),
    .io_co(FullAdder_33_io_co)
  );
  FullAdder FullAdder_34 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_34_io_a),
    .io_b(FullAdder_34_io_b),
    .io_ci(FullAdder_34_io_ci),
    .io_s(FullAdder_34_io_s),
    .io_co(FullAdder_34_io_co)
  );
  FullAdder FullAdder_35 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_35_io_a),
    .io_b(FullAdder_35_io_b),
    .io_ci(FullAdder_35_io_ci),
    .io_s(FullAdder_35_io_s),
    .io_co(FullAdder_35_io_co)
  );
  FullAdder FullAdder_36 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_36_io_a),
    .io_b(FullAdder_36_io_b),
    .io_ci(FullAdder_36_io_ci),
    .io_s(FullAdder_36_io_s),
    .io_co(FullAdder_36_io_co)
  );
  FullAdder FullAdder_37 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_37_io_a),
    .io_b(FullAdder_37_io_b),
    .io_ci(FullAdder_37_io_ci),
    .io_s(FullAdder_37_io_s),
    .io_co(FullAdder_37_io_co)
  );
  FullAdder FullAdder_38 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_38_io_a),
    .io_b(FullAdder_38_io_b),
    .io_ci(FullAdder_38_io_ci),
    .io_s(FullAdder_38_io_s),
    .io_co(FullAdder_38_io_co)
  );
  FullAdder FullAdder_39 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_39_io_a),
    .io_b(FullAdder_39_io_b),
    .io_ci(FullAdder_39_io_ci),
    .io_s(FullAdder_39_io_s),
    .io_co(FullAdder_39_io_co)
  );
  FullAdder FullAdder_40 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_40_io_a),
    .io_b(FullAdder_40_io_b),
    .io_ci(FullAdder_40_io_ci),
    .io_s(FullAdder_40_io_s),
    .io_co(FullAdder_40_io_co)
  );
  FullAdder FullAdder_41 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_41_io_a),
    .io_b(FullAdder_41_io_b),
    .io_ci(FullAdder_41_io_ci),
    .io_s(FullAdder_41_io_s),
    .io_co(FullAdder_41_io_co)
  );
  FullAdder FullAdder_42 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_42_io_a),
    .io_b(FullAdder_42_io_b),
    .io_ci(FullAdder_42_io_ci),
    .io_s(FullAdder_42_io_s),
    .io_co(FullAdder_42_io_co)
  );
  FullAdder FullAdder_43 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_43_io_a),
    .io_b(FullAdder_43_io_b),
    .io_ci(FullAdder_43_io_ci),
    .io_s(FullAdder_43_io_s),
    .io_co(FullAdder_43_io_co)
  );
  FullAdder FullAdder_44 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_44_io_a),
    .io_b(FullAdder_44_io_b),
    .io_ci(FullAdder_44_io_ci),
    .io_s(FullAdder_44_io_s),
    .io_co(FullAdder_44_io_co)
  );
  FullAdder FullAdder_45 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_45_io_a),
    .io_b(FullAdder_45_io_b),
    .io_ci(FullAdder_45_io_ci),
    .io_s(FullAdder_45_io_s),
    .io_co(FullAdder_45_io_co)
  );
  FullAdder FullAdder_46 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_46_io_a),
    .io_b(FullAdder_46_io_b),
    .io_ci(FullAdder_46_io_ci),
    .io_s(FullAdder_46_io_s),
    .io_co(FullAdder_46_io_co)
  );
  FullAdder FullAdder_47 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_47_io_a),
    .io_b(FullAdder_47_io_b),
    .io_ci(FullAdder_47_io_ci),
    .io_s(FullAdder_47_io_s),
    .io_co(FullAdder_47_io_co)
  );
  FullAdder FullAdder_48 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_48_io_a),
    .io_b(FullAdder_48_io_b),
    .io_ci(FullAdder_48_io_ci),
    .io_s(FullAdder_48_io_s),
    .io_co(FullAdder_48_io_co)
  );
  FullAdder FullAdder_49 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_49_io_a),
    .io_b(FullAdder_49_io_b),
    .io_ci(FullAdder_49_io_ci),
    .io_s(FullAdder_49_io_s),
    .io_co(FullAdder_49_io_co)
  );
  FullAdder FullAdder_50 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_50_io_a),
    .io_b(FullAdder_50_io_b),
    .io_ci(FullAdder_50_io_ci),
    .io_s(FullAdder_50_io_s),
    .io_co(FullAdder_50_io_co)
  );
  FullAdder FullAdder_51 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_51_io_a),
    .io_b(FullAdder_51_io_b),
    .io_ci(FullAdder_51_io_ci),
    .io_s(FullAdder_51_io_s),
    .io_co(FullAdder_51_io_co)
  );
  FullAdder FullAdder_52 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_52_io_a),
    .io_b(FullAdder_52_io_b),
    .io_ci(FullAdder_52_io_ci),
    .io_s(FullAdder_52_io_s),
    .io_co(FullAdder_52_io_co)
  );
  FullAdder FullAdder_53 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_53_io_a),
    .io_b(FullAdder_53_io_b),
    .io_ci(FullAdder_53_io_ci),
    .io_s(FullAdder_53_io_s),
    .io_co(FullAdder_53_io_co)
  );
  FullAdder FullAdder_54 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_54_io_a),
    .io_b(FullAdder_54_io_b),
    .io_ci(FullAdder_54_io_ci),
    .io_s(FullAdder_54_io_s),
    .io_co(FullAdder_54_io_co)
  );
  FullAdder FullAdder_55 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_55_io_a),
    .io_b(FullAdder_55_io_b),
    .io_ci(FullAdder_55_io_ci),
    .io_s(FullAdder_55_io_s),
    .io_co(FullAdder_55_io_co)
  );
  FullAdder FullAdder_56 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_56_io_a),
    .io_b(FullAdder_56_io_b),
    .io_ci(FullAdder_56_io_ci),
    .io_s(FullAdder_56_io_s),
    .io_co(FullAdder_56_io_co)
  );
  FullAdder FullAdder_57 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_57_io_a),
    .io_b(FullAdder_57_io_b),
    .io_ci(FullAdder_57_io_ci),
    .io_s(FullAdder_57_io_s),
    .io_co(FullAdder_57_io_co)
  );
  FullAdder FullAdder_58 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_58_io_a),
    .io_b(FullAdder_58_io_b),
    .io_ci(FullAdder_58_io_ci),
    .io_s(FullAdder_58_io_s),
    .io_co(FullAdder_58_io_co)
  );
  FullAdder FullAdder_59 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_59_io_a),
    .io_b(FullAdder_59_io_b),
    .io_ci(FullAdder_59_io_ci),
    .io_s(FullAdder_59_io_s),
    .io_co(FullAdder_59_io_co)
  );
  FullAdder FullAdder_60 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_60_io_a),
    .io_b(FullAdder_60_io_b),
    .io_ci(FullAdder_60_io_ci),
    .io_s(FullAdder_60_io_s),
    .io_co(FullAdder_60_io_co)
  );
  FullAdder FullAdder_61 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_61_io_a),
    .io_b(FullAdder_61_io_b),
    .io_ci(FullAdder_61_io_ci),
    .io_s(FullAdder_61_io_s),
    .io_co(FullAdder_61_io_co)
  );
  FullAdder FullAdder_62 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_62_io_a),
    .io_b(FullAdder_62_io_b),
    .io_ci(FullAdder_62_io_ci),
    .io_s(FullAdder_62_io_s),
    .io_co(FullAdder_62_io_co)
  );
  FullAdder FullAdder_63 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_63_io_a),
    .io_b(FullAdder_63_io_b),
    .io_ci(FullAdder_63_io_ci),
    .io_s(FullAdder_63_io_s),
    .io_co(FullAdder_63_io_co)
  );
  FullAdder FullAdder_64 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_64_io_a),
    .io_b(FullAdder_64_io_b),
    .io_ci(FullAdder_64_io_ci),
    .io_s(FullAdder_64_io_s),
    .io_co(FullAdder_64_io_co)
  );
  FullAdder FullAdder_65 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_65_io_a),
    .io_b(FullAdder_65_io_b),
    .io_ci(FullAdder_65_io_ci),
    .io_s(FullAdder_65_io_s),
    .io_co(FullAdder_65_io_co)
  );
  FullAdder FullAdder_66 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_66_io_a),
    .io_b(FullAdder_66_io_b),
    .io_ci(FullAdder_66_io_ci),
    .io_s(FullAdder_66_io_s),
    .io_co(FullAdder_66_io_co)
  );
  FullAdder FullAdder_67 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_67_io_a),
    .io_b(FullAdder_67_io_b),
    .io_ci(FullAdder_67_io_ci),
    .io_s(FullAdder_67_io_s),
    .io_co(FullAdder_67_io_co)
  );
  FullAdder FullAdder_68 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_68_io_a),
    .io_b(FullAdder_68_io_b),
    .io_ci(FullAdder_68_io_ci),
    .io_s(FullAdder_68_io_s),
    .io_co(FullAdder_68_io_co)
  );
  FullAdder FullAdder_69 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_69_io_a),
    .io_b(FullAdder_69_io_b),
    .io_ci(FullAdder_69_io_ci),
    .io_s(FullAdder_69_io_s),
    .io_co(FullAdder_69_io_co)
  );
  FullAdder FullAdder_70 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_70_io_a),
    .io_b(FullAdder_70_io_b),
    .io_ci(FullAdder_70_io_ci),
    .io_s(FullAdder_70_io_s),
    .io_co(FullAdder_70_io_co)
  );
  FullAdder FullAdder_71 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_71_io_a),
    .io_b(FullAdder_71_io_b),
    .io_ci(FullAdder_71_io_ci),
    .io_s(FullAdder_71_io_s),
    .io_co(FullAdder_71_io_co)
  );
  FullAdder FullAdder_72 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_72_io_a),
    .io_b(FullAdder_72_io_b),
    .io_ci(FullAdder_72_io_ci),
    .io_s(FullAdder_72_io_s),
    .io_co(FullAdder_72_io_co)
  );
  FullAdder FullAdder_73 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_73_io_a),
    .io_b(FullAdder_73_io_b),
    .io_ci(FullAdder_73_io_ci),
    .io_s(FullAdder_73_io_s),
    .io_co(FullAdder_73_io_co)
  );
  FullAdder FullAdder_74 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_74_io_a),
    .io_b(FullAdder_74_io_b),
    .io_ci(FullAdder_74_io_ci),
    .io_s(FullAdder_74_io_s),
    .io_co(FullAdder_74_io_co)
  );
  FullAdder FullAdder_75 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_75_io_a),
    .io_b(FullAdder_75_io_b),
    .io_ci(FullAdder_75_io_ci),
    .io_s(FullAdder_75_io_s),
    .io_co(FullAdder_75_io_co)
  );
  FullAdder FullAdder_76 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_76_io_a),
    .io_b(FullAdder_76_io_b),
    .io_ci(FullAdder_76_io_ci),
    .io_s(FullAdder_76_io_s),
    .io_co(FullAdder_76_io_co)
  );
  FullAdder FullAdder_77 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_77_io_a),
    .io_b(FullAdder_77_io_b),
    .io_ci(FullAdder_77_io_ci),
    .io_s(FullAdder_77_io_s),
    .io_co(FullAdder_77_io_co)
  );
  FullAdder FullAdder_78 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_78_io_a),
    .io_b(FullAdder_78_io_b),
    .io_ci(FullAdder_78_io_ci),
    .io_s(FullAdder_78_io_s),
    .io_co(FullAdder_78_io_co)
  );
  FullAdder FullAdder_79 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_79_io_a),
    .io_b(FullAdder_79_io_b),
    .io_ci(FullAdder_79_io_ci),
    .io_s(FullAdder_79_io_s),
    .io_co(FullAdder_79_io_co)
  );
  FullAdder FullAdder_80 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_80_io_a),
    .io_b(FullAdder_80_io_b),
    .io_ci(FullAdder_80_io_ci),
    .io_s(FullAdder_80_io_s),
    .io_co(FullAdder_80_io_co)
  );
  FullAdder FullAdder_81 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_81_io_a),
    .io_b(FullAdder_81_io_b),
    .io_ci(FullAdder_81_io_ci),
    .io_s(FullAdder_81_io_s),
    .io_co(FullAdder_81_io_co)
  );
  FullAdder FullAdder_82 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_82_io_a),
    .io_b(FullAdder_82_io_b),
    .io_ci(FullAdder_82_io_ci),
    .io_s(FullAdder_82_io_s),
    .io_co(FullAdder_82_io_co)
  );
  FullAdder FullAdder_83 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_83_io_a),
    .io_b(FullAdder_83_io_b),
    .io_ci(FullAdder_83_io_ci),
    .io_s(FullAdder_83_io_s),
    .io_co(FullAdder_83_io_co)
  );
  FullAdder FullAdder_84 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_84_io_a),
    .io_b(FullAdder_84_io_b),
    .io_ci(FullAdder_84_io_ci),
    .io_s(FullAdder_84_io_s),
    .io_co(FullAdder_84_io_co)
  );
  FullAdder FullAdder_85 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_85_io_a),
    .io_b(FullAdder_85_io_b),
    .io_ci(FullAdder_85_io_ci),
    .io_s(FullAdder_85_io_s),
    .io_co(FullAdder_85_io_co)
  );
  FullAdder FullAdder_86 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_86_io_a),
    .io_b(FullAdder_86_io_b),
    .io_ci(FullAdder_86_io_ci),
    .io_s(FullAdder_86_io_s),
    .io_co(FullAdder_86_io_co)
  );
  FullAdder FullAdder_87 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_87_io_a),
    .io_b(FullAdder_87_io_b),
    .io_ci(FullAdder_87_io_ci),
    .io_s(FullAdder_87_io_s),
    .io_co(FullAdder_87_io_co)
  );
  FullAdder FullAdder_88 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_88_io_a),
    .io_b(FullAdder_88_io_b),
    .io_ci(FullAdder_88_io_ci),
    .io_s(FullAdder_88_io_s),
    .io_co(FullAdder_88_io_co)
  );
  FullAdder FullAdder_89 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_89_io_a),
    .io_b(FullAdder_89_io_b),
    .io_ci(FullAdder_89_io_ci),
    .io_s(FullAdder_89_io_s),
    .io_co(FullAdder_89_io_co)
  );
  FullAdder FullAdder_90 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_90_io_a),
    .io_b(FullAdder_90_io_b),
    .io_ci(FullAdder_90_io_ci),
    .io_s(FullAdder_90_io_s),
    .io_co(FullAdder_90_io_co)
  );
  FullAdder FullAdder_91 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_91_io_a),
    .io_b(FullAdder_91_io_b),
    .io_ci(FullAdder_91_io_ci),
    .io_s(FullAdder_91_io_s),
    .io_co(FullAdder_91_io_co)
  );
  FullAdder FullAdder_92 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_92_io_a),
    .io_b(FullAdder_92_io_b),
    .io_ci(FullAdder_92_io_ci),
    .io_s(FullAdder_92_io_s),
    .io_co(FullAdder_92_io_co)
  );
  FullAdder FullAdder_93 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_93_io_a),
    .io_b(FullAdder_93_io_b),
    .io_ci(FullAdder_93_io_ci),
    .io_s(FullAdder_93_io_s),
    .io_co(FullAdder_93_io_co)
  );
  FullAdder FullAdder_94 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_94_io_a),
    .io_b(FullAdder_94_io_b),
    .io_ci(FullAdder_94_io_ci),
    .io_s(FullAdder_94_io_s),
    .io_co(FullAdder_94_io_co)
  );
  FullAdder FullAdder_95 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_95_io_a),
    .io_b(FullAdder_95_io_b),
    .io_ci(FullAdder_95_io_ci),
    .io_s(FullAdder_95_io_s),
    .io_co(FullAdder_95_io_co)
  );
  FullAdder FullAdder_96 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_96_io_a),
    .io_b(FullAdder_96_io_b),
    .io_ci(FullAdder_96_io_ci),
    .io_s(FullAdder_96_io_s),
    .io_co(FullAdder_96_io_co)
  );
  FullAdder FullAdder_97 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_97_io_a),
    .io_b(FullAdder_97_io_b),
    .io_ci(FullAdder_97_io_ci),
    .io_s(FullAdder_97_io_s),
    .io_co(FullAdder_97_io_co)
  );
  FullAdder FullAdder_98 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_98_io_a),
    .io_b(FullAdder_98_io_b),
    .io_ci(FullAdder_98_io_ci),
    .io_s(FullAdder_98_io_s),
    .io_co(FullAdder_98_io_co)
  );
  FullAdder FullAdder_99 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_99_io_a),
    .io_b(FullAdder_99_io_b),
    .io_ci(FullAdder_99_io_ci),
    .io_s(FullAdder_99_io_s),
    .io_co(FullAdder_99_io_co)
  );
  FullAdder FullAdder_100 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_100_io_a),
    .io_b(FullAdder_100_io_b),
    .io_ci(FullAdder_100_io_ci),
    .io_s(FullAdder_100_io_s),
    .io_co(FullAdder_100_io_co)
  );
  FullAdder FullAdder_101 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_101_io_a),
    .io_b(FullAdder_101_io_b),
    .io_ci(FullAdder_101_io_ci),
    .io_s(FullAdder_101_io_s),
    .io_co(FullAdder_101_io_co)
  );
  FullAdder FullAdder_102 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_102_io_a),
    .io_b(FullAdder_102_io_b),
    .io_ci(FullAdder_102_io_ci),
    .io_s(FullAdder_102_io_s),
    .io_co(FullAdder_102_io_co)
  );
  FullAdder FullAdder_103 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_103_io_a),
    .io_b(FullAdder_103_io_b),
    .io_ci(FullAdder_103_io_ci),
    .io_s(FullAdder_103_io_s),
    .io_co(FullAdder_103_io_co)
  );
  FullAdder FullAdder_104 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_104_io_a),
    .io_b(FullAdder_104_io_b),
    .io_ci(FullAdder_104_io_ci),
    .io_s(FullAdder_104_io_s),
    .io_co(FullAdder_104_io_co)
  );
  FullAdder FullAdder_105 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_105_io_a),
    .io_b(FullAdder_105_io_b),
    .io_ci(FullAdder_105_io_ci),
    .io_s(FullAdder_105_io_s),
    .io_co(FullAdder_105_io_co)
  );
  FullAdder FullAdder_106 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_106_io_a),
    .io_b(FullAdder_106_io_b),
    .io_ci(FullAdder_106_io_ci),
    .io_s(FullAdder_106_io_s),
    .io_co(FullAdder_106_io_co)
  );
  FullAdder FullAdder_107 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_107_io_a),
    .io_b(FullAdder_107_io_b),
    .io_ci(FullAdder_107_io_ci),
    .io_s(FullAdder_107_io_s),
    .io_co(FullAdder_107_io_co)
  );
  FullAdder FullAdder_108 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_108_io_a),
    .io_b(FullAdder_108_io_b),
    .io_ci(FullAdder_108_io_ci),
    .io_s(FullAdder_108_io_s),
    .io_co(FullAdder_108_io_co)
  );
  FullAdder FullAdder_109 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_109_io_a),
    .io_b(FullAdder_109_io_b),
    .io_ci(FullAdder_109_io_ci),
    .io_s(FullAdder_109_io_s),
    .io_co(FullAdder_109_io_co)
  );
  FullAdder FullAdder_110 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_110_io_a),
    .io_b(FullAdder_110_io_b),
    .io_ci(FullAdder_110_io_ci),
    .io_s(FullAdder_110_io_s),
    .io_co(FullAdder_110_io_co)
  );
  FullAdder FullAdder_111 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_111_io_a),
    .io_b(FullAdder_111_io_b),
    .io_ci(FullAdder_111_io_ci),
    .io_s(FullAdder_111_io_s),
    .io_co(FullAdder_111_io_co)
  );
  FullAdder FullAdder_112 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_112_io_a),
    .io_b(FullAdder_112_io_b),
    .io_ci(FullAdder_112_io_ci),
    .io_s(FullAdder_112_io_s),
    .io_co(FullAdder_112_io_co)
  );
  FullAdder FullAdder_113 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_113_io_a),
    .io_b(FullAdder_113_io_b),
    .io_ci(FullAdder_113_io_ci),
    .io_s(FullAdder_113_io_s),
    .io_co(FullAdder_113_io_co)
  );
  FullAdder FullAdder_114 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_114_io_a),
    .io_b(FullAdder_114_io_b),
    .io_ci(FullAdder_114_io_ci),
    .io_s(FullAdder_114_io_s),
    .io_co(FullAdder_114_io_co)
  );
  FullAdder FullAdder_115 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_115_io_a),
    .io_b(FullAdder_115_io_b),
    .io_ci(FullAdder_115_io_ci),
    .io_s(FullAdder_115_io_s),
    .io_co(FullAdder_115_io_co)
  );
  FullAdder FullAdder_116 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_116_io_a),
    .io_b(FullAdder_116_io_b),
    .io_ci(FullAdder_116_io_ci),
    .io_s(FullAdder_116_io_s),
    .io_co(FullAdder_116_io_co)
  );
  FullAdder FullAdder_117 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_117_io_a),
    .io_b(FullAdder_117_io_b),
    .io_ci(FullAdder_117_io_ci),
    .io_s(FullAdder_117_io_s),
    .io_co(FullAdder_117_io_co)
  );
  FullAdder FullAdder_118 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_118_io_a),
    .io_b(FullAdder_118_io_b),
    .io_ci(FullAdder_118_io_ci),
    .io_s(FullAdder_118_io_s),
    .io_co(FullAdder_118_io_co)
  );
  FullAdder FullAdder_119 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_119_io_a),
    .io_b(FullAdder_119_io_b),
    .io_ci(FullAdder_119_io_ci),
    .io_s(FullAdder_119_io_s),
    .io_co(FullAdder_119_io_co)
  );
  FullAdder FullAdder_120 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_120_io_a),
    .io_b(FullAdder_120_io_b),
    .io_ci(FullAdder_120_io_ci),
    .io_s(FullAdder_120_io_s),
    .io_co(FullAdder_120_io_co)
  );
  FullAdder FullAdder_121 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_121_io_a),
    .io_b(FullAdder_121_io_b),
    .io_ci(FullAdder_121_io_ci),
    .io_s(FullAdder_121_io_s),
    .io_co(FullAdder_121_io_co)
  );
  FullAdder FullAdder_122 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_122_io_a),
    .io_b(FullAdder_122_io_b),
    .io_ci(FullAdder_122_io_ci),
    .io_s(FullAdder_122_io_s),
    .io_co(FullAdder_122_io_co)
  );
  FullAdder FullAdder_123 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_123_io_a),
    .io_b(FullAdder_123_io_b),
    .io_ci(FullAdder_123_io_ci),
    .io_s(FullAdder_123_io_s),
    .io_co(FullAdder_123_io_co)
  );
  FullAdder FullAdder_124 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_124_io_a),
    .io_b(FullAdder_124_io_b),
    .io_ci(FullAdder_124_io_ci),
    .io_s(FullAdder_124_io_s),
    .io_co(FullAdder_124_io_co)
  );
  FullAdder FullAdder_125 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_125_io_a),
    .io_b(FullAdder_125_io_b),
    .io_ci(FullAdder_125_io_ci),
    .io_s(FullAdder_125_io_s),
    .io_co(FullAdder_125_io_co)
  );
  FullAdder FullAdder_126 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_126_io_a),
    .io_b(FullAdder_126_io_b),
    .io_ci(FullAdder_126_io_ci),
    .io_s(FullAdder_126_io_s),
    .io_co(FullAdder_126_io_co)
  );
  FullAdder FullAdder_127 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_127_io_a),
    .io_b(FullAdder_127_io_b),
    .io_ci(FullAdder_127_io_ci),
    .io_s(FullAdder_127_io_s),
    .io_co(FullAdder_127_io_co)
  );
  FullAdder FullAdder_128 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_128_io_a),
    .io_b(FullAdder_128_io_b),
    .io_ci(FullAdder_128_io_ci),
    .io_s(FullAdder_128_io_s),
    .io_co(FullAdder_128_io_co)
  );
  FullAdder FullAdder_129 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_129_io_a),
    .io_b(FullAdder_129_io_b),
    .io_ci(FullAdder_129_io_ci),
    .io_s(FullAdder_129_io_s),
    .io_co(FullAdder_129_io_co)
  );
  FullAdder FullAdder_130 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_130_io_a),
    .io_b(FullAdder_130_io_b),
    .io_ci(FullAdder_130_io_ci),
    .io_s(FullAdder_130_io_s),
    .io_co(FullAdder_130_io_co)
  );
  FullAdder FullAdder_131 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_131_io_a),
    .io_b(FullAdder_131_io_b),
    .io_ci(FullAdder_131_io_ci),
    .io_s(FullAdder_131_io_s),
    .io_co(FullAdder_131_io_co)
  );
  FullAdder FullAdder_132 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_132_io_a),
    .io_b(FullAdder_132_io_b),
    .io_ci(FullAdder_132_io_ci),
    .io_s(FullAdder_132_io_s),
    .io_co(FullAdder_132_io_co)
  );
  FullAdder FullAdder_133 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_133_io_a),
    .io_b(FullAdder_133_io_b),
    .io_ci(FullAdder_133_io_ci),
    .io_s(FullAdder_133_io_s),
    .io_co(FullAdder_133_io_co)
  );
  FullAdder FullAdder_134 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_134_io_a),
    .io_b(FullAdder_134_io_b),
    .io_ci(FullAdder_134_io_ci),
    .io_s(FullAdder_134_io_s),
    .io_co(FullAdder_134_io_co)
  );
  FullAdder FullAdder_135 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_135_io_a),
    .io_b(FullAdder_135_io_b),
    .io_ci(FullAdder_135_io_ci),
    .io_s(FullAdder_135_io_s),
    .io_co(FullAdder_135_io_co)
  );
  FullAdder FullAdder_136 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_136_io_a),
    .io_b(FullAdder_136_io_b),
    .io_ci(FullAdder_136_io_ci),
    .io_s(FullAdder_136_io_s),
    .io_co(FullAdder_136_io_co)
  );
  FullAdder FullAdder_137 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_137_io_a),
    .io_b(FullAdder_137_io_b),
    .io_ci(FullAdder_137_io_ci),
    .io_s(FullAdder_137_io_s),
    .io_co(FullAdder_137_io_co)
  );
  FullAdder FullAdder_138 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_138_io_a),
    .io_b(FullAdder_138_io_b),
    .io_ci(FullAdder_138_io_ci),
    .io_s(FullAdder_138_io_s),
    .io_co(FullAdder_138_io_co)
  );
  FullAdder FullAdder_139 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_139_io_a),
    .io_b(FullAdder_139_io_b),
    .io_ci(FullAdder_139_io_ci),
    .io_s(FullAdder_139_io_s),
    .io_co(FullAdder_139_io_co)
  );
  FullAdder FullAdder_140 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_140_io_a),
    .io_b(FullAdder_140_io_b),
    .io_ci(FullAdder_140_io_ci),
    .io_s(FullAdder_140_io_s),
    .io_co(FullAdder_140_io_co)
  );
  FullAdder FullAdder_141 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_141_io_a),
    .io_b(FullAdder_141_io_b),
    .io_ci(FullAdder_141_io_ci),
    .io_s(FullAdder_141_io_s),
    .io_co(FullAdder_141_io_co)
  );
  FullAdder FullAdder_142 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_142_io_a),
    .io_b(FullAdder_142_io_b),
    .io_ci(FullAdder_142_io_ci),
    .io_s(FullAdder_142_io_s),
    .io_co(FullAdder_142_io_co)
  );
  FullAdder FullAdder_143 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_143_io_a),
    .io_b(FullAdder_143_io_b),
    .io_ci(FullAdder_143_io_ci),
    .io_s(FullAdder_143_io_s),
    .io_co(FullAdder_143_io_co)
  );
  FullAdder FullAdder_144 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_144_io_a),
    .io_b(FullAdder_144_io_b),
    .io_ci(FullAdder_144_io_ci),
    .io_s(FullAdder_144_io_s),
    .io_co(FullAdder_144_io_co)
  );
  FullAdder FullAdder_145 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_145_io_a),
    .io_b(FullAdder_145_io_b),
    .io_ci(FullAdder_145_io_ci),
    .io_s(FullAdder_145_io_s),
    .io_co(FullAdder_145_io_co)
  );
  FullAdder FullAdder_146 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_146_io_a),
    .io_b(FullAdder_146_io_b),
    .io_ci(FullAdder_146_io_ci),
    .io_s(FullAdder_146_io_s),
    .io_co(FullAdder_146_io_co)
  );
  FullAdder FullAdder_147 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_147_io_a),
    .io_b(FullAdder_147_io_b),
    .io_ci(FullAdder_147_io_ci),
    .io_s(FullAdder_147_io_s),
    .io_co(FullAdder_147_io_co)
  );
  FullAdder FullAdder_148 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_148_io_a),
    .io_b(FullAdder_148_io_b),
    .io_ci(FullAdder_148_io_ci),
    .io_s(FullAdder_148_io_s),
    .io_co(FullAdder_148_io_co)
  );
  FullAdder FullAdder_149 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_149_io_a),
    .io_b(FullAdder_149_io_b),
    .io_ci(FullAdder_149_io_ci),
    .io_s(FullAdder_149_io_s),
    .io_co(FullAdder_149_io_co)
  );
  FullAdder FullAdder_150 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_150_io_a),
    .io_b(FullAdder_150_io_b),
    .io_ci(FullAdder_150_io_ci),
    .io_s(FullAdder_150_io_s),
    .io_co(FullAdder_150_io_co)
  );
  FullAdder FullAdder_151 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_151_io_a),
    .io_b(FullAdder_151_io_b),
    .io_ci(FullAdder_151_io_ci),
    .io_s(FullAdder_151_io_s),
    .io_co(FullAdder_151_io_co)
  );
  FullAdder FullAdder_152 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_152_io_a),
    .io_b(FullAdder_152_io_b),
    .io_ci(FullAdder_152_io_ci),
    .io_s(FullAdder_152_io_s),
    .io_co(FullAdder_152_io_co)
  );
  FullAdder FullAdder_153 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_153_io_a),
    .io_b(FullAdder_153_io_b),
    .io_ci(FullAdder_153_io_ci),
    .io_s(FullAdder_153_io_s),
    .io_co(FullAdder_153_io_co)
  );
  HalfAdder HalfAdder ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_io_a),
    .io_b(HalfAdder_io_b),
    .io_s(HalfAdder_io_s),
    .io_co(HalfAdder_io_co)
  );
  FullAdder FullAdder_154 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_154_io_a),
    .io_b(FullAdder_154_io_b),
    .io_ci(FullAdder_154_io_ci),
    .io_s(FullAdder_154_io_s),
    .io_co(FullAdder_154_io_co)
  );
  FullAdder FullAdder_155 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_155_io_a),
    .io_b(FullAdder_155_io_b),
    .io_ci(FullAdder_155_io_ci),
    .io_s(FullAdder_155_io_s),
    .io_co(FullAdder_155_io_co)
  );
  FullAdder FullAdder_156 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_156_io_a),
    .io_b(FullAdder_156_io_b),
    .io_ci(FullAdder_156_io_ci),
    .io_s(FullAdder_156_io_s),
    .io_co(FullAdder_156_io_co)
  );
  FullAdder FullAdder_157 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_157_io_a),
    .io_b(FullAdder_157_io_b),
    .io_ci(FullAdder_157_io_ci),
    .io_s(FullAdder_157_io_s),
    .io_co(FullAdder_157_io_co)
  );
  FullAdder FullAdder_158 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_158_io_a),
    .io_b(FullAdder_158_io_b),
    .io_ci(FullAdder_158_io_ci),
    .io_s(FullAdder_158_io_s),
    .io_co(FullAdder_158_io_co)
  );
  FullAdder FullAdder_159 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_159_io_a),
    .io_b(FullAdder_159_io_b),
    .io_ci(FullAdder_159_io_ci),
    .io_s(FullAdder_159_io_s),
    .io_co(FullAdder_159_io_co)
  );
  FullAdder FullAdder_160 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_160_io_a),
    .io_b(FullAdder_160_io_b),
    .io_ci(FullAdder_160_io_ci),
    .io_s(FullAdder_160_io_s),
    .io_co(FullAdder_160_io_co)
  );
  FullAdder FullAdder_161 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_161_io_a),
    .io_b(FullAdder_161_io_b),
    .io_ci(FullAdder_161_io_ci),
    .io_s(FullAdder_161_io_s),
    .io_co(FullAdder_161_io_co)
  );
  FullAdder FullAdder_162 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_162_io_a),
    .io_b(FullAdder_162_io_b),
    .io_ci(FullAdder_162_io_ci),
    .io_s(FullAdder_162_io_s),
    .io_co(FullAdder_162_io_co)
  );
  FullAdder FullAdder_163 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_163_io_a),
    .io_b(FullAdder_163_io_b),
    .io_ci(FullAdder_163_io_ci),
    .io_s(FullAdder_163_io_s),
    .io_co(FullAdder_163_io_co)
  );
  FullAdder FullAdder_164 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_164_io_a),
    .io_b(FullAdder_164_io_b),
    .io_ci(FullAdder_164_io_ci),
    .io_s(FullAdder_164_io_s),
    .io_co(FullAdder_164_io_co)
  );
  FullAdder FullAdder_165 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_165_io_a),
    .io_b(FullAdder_165_io_b),
    .io_ci(FullAdder_165_io_ci),
    .io_s(FullAdder_165_io_s),
    .io_co(FullAdder_165_io_co)
  );
  FullAdder FullAdder_166 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_166_io_a),
    .io_b(FullAdder_166_io_b),
    .io_ci(FullAdder_166_io_ci),
    .io_s(FullAdder_166_io_s),
    .io_co(FullAdder_166_io_co)
  );
  FullAdder FullAdder_167 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_167_io_a),
    .io_b(FullAdder_167_io_b),
    .io_ci(FullAdder_167_io_ci),
    .io_s(FullAdder_167_io_s),
    .io_co(FullAdder_167_io_co)
  );
  FullAdder FullAdder_168 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_168_io_a),
    .io_b(FullAdder_168_io_b),
    .io_ci(FullAdder_168_io_ci),
    .io_s(FullAdder_168_io_s),
    .io_co(FullAdder_168_io_co)
  );
  FullAdder FullAdder_169 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_169_io_a),
    .io_b(FullAdder_169_io_b),
    .io_ci(FullAdder_169_io_ci),
    .io_s(FullAdder_169_io_s),
    .io_co(FullAdder_169_io_co)
  );
  FullAdder FullAdder_170 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_170_io_a),
    .io_b(FullAdder_170_io_b),
    .io_ci(FullAdder_170_io_ci),
    .io_s(FullAdder_170_io_s),
    .io_co(FullAdder_170_io_co)
  );
  FullAdder FullAdder_171 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_171_io_a),
    .io_b(FullAdder_171_io_b),
    .io_ci(FullAdder_171_io_ci),
    .io_s(FullAdder_171_io_s),
    .io_co(FullAdder_171_io_co)
  );
  FullAdder FullAdder_172 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_172_io_a),
    .io_b(FullAdder_172_io_b),
    .io_ci(FullAdder_172_io_ci),
    .io_s(FullAdder_172_io_s),
    .io_co(FullAdder_172_io_co)
  );
  FullAdder FullAdder_173 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_173_io_a),
    .io_b(FullAdder_173_io_b),
    .io_ci(FullAdder_173_io_ci),
    .io_s(FullAdder_173_io_s),
    .io_co(FullAdder_173_io_co)
  );
  FullAdder FullAdder_174 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_174_io_a),
    .io_b(FullAdder_174_io_b),
    .io_ci(FullAdder_174_io_ci),
    .io_s(FullAdder_174_io_s),
    .io_co(FullAdder_174_io_co)
  );
  HalfAdder HalfAdder_1 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_1_io_a),
    .io_b(HalfAdder_1_io_b),
    .io_s(HalfAdder_1_io_s),
    .io_co(HalfAdder_1_io_co)
  );
  FullAdder FullAdder_175 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_175_io_a),
    .io_b(FullAdder_175_io_b),
    .io_ci(FullAdder_175_io_ci),
    .io_s(FullAdder_175_io_s),
    .io_co(FullAdder_175_io_co)
  );
  FullAdder FullAdder_176 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_176_io_a),
    .io_b(FullAdder_176_io_b),
    .io_ci(FullAdder_176_io_ci),
    .io_s(FullAdder_176_io_s),
    .io_co(FullAdder_176_io_co)
  );
  FullAdder FullAdder_177 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_177_io_a),
    .io_b(FullAdder_177_io_b),
    .io_ci(FullAdder_177_io_ci),
    .io_s(FullAdder_177_io_s),
    .io_co(FullAdder_177_io_co)
  );
  FullAdder FullAdder_178 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_178_io_a),
    .io_b(FullAdder_178_io_b),
    .io_ci(FullAdder_178_io_ci),
    .io_s(FullAdder_178_io_s),
    .io_co(FullAdder_178_io_co)
  );
  FullAdder FullAdder_179 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_179_io_a),
    .io_b(FullAdder_179_io_b),
    .io_ci(FullAdder_179_io_ci),
    .io_s(FullAdder_179_io_s),
    .io_co(FullAdder_179_io_co)
  );
  FullAdder FullAdder_180 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_180_io_a),
    .io_b(FullAdder_180_io_b),
    .io_ci(FullAdder_180_io_ci),
    .io_s(FullAdder_180_io_s),
    .io_co(FullAdder_180_io_co)
  );
  FullAdder FullAdder_181 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_181_io_a),
    .io_b(FullAdder_181_io_b),
    .io_ci(FullAdder_181_io_ci),
    .io_s(FullAdder_181_io_s),
    .io_co(FullAdder_181_io_co)
  );
  FullAdder FullAdder_182 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_182_io_a),
    .io_b(FullAdder_182_io_b),
    .io_ci(FullAdder_182_io_ci),
    .io_s(FullAdder_182_io_s),
    .io_co(FullAdder_182_io_co)
  );
  FullAdder FullAdder_183 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_183_io_a),
    .io_b(FullAdder_183_io_b),
    .io_ci(FullAdder_183_io_ci),
    .io_s(FullAdder_183_io_s),
    .io_co(FullAdder_183_io_co)
  );
  FullAdder FullAdder_184 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_184_io_a),
    .io_b(FullAdder_184_io_b),
    .io_ci(FullAdder_184_io_ci),
    .io_s(FullAdder_184_io_s),
    .io_co(FullAdder_184_io_co)
  );
  FullAdder FullAdder_185 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_185_io_a),
    .io_b(FullAdder_185_io_b),
    .io_ci(FullAdder_185_io_ci),
    .io_s(FullAdder_185_io_s),
    .io_co(FullAdder_185_io_co)
  );
  FullAdder FullAdder_186 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_186_io_a),
    .io_b(FullAdder_186_io_b),
    .io_ci(FullAdder_186_io_ci),
    .io_s(FullAdder_186_io_s),
    .io_co(FullAdder_186_io_co)
  );
  FullAdder FullAdder_187 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_187_io_a),
    .io_b(FullAdder_187_io_b),
    .io_ci(FullAdder_187_io_ci),
    .io_s(FullAdder_187_io_s),
    .io_co(FullAdder_187_io_co)
  );
  HalfAdder HalfAdder_2 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_2_io_a),
    .io_b(HalfAdder_2_io_b),
    .io_s(HalfAdder_2_io_s),
    .io_co(HalfAdder_2_io_co)
  );
  FullAdder FullAdder_188 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_188_io_a),
    .io_b(FullAdder_188_io_b),
    .io_ci(FullAdder_188_io_ci),
    .io_s(FullAdder_188_io_s),
    .io_co(FullAdder_188_io_co)
  );
  FullAdder FullAdder_189 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_189_io_a),
    .io_b(FullAdder_189_io_b),
    .io_ci(FullAdder_189_io_ci),
    .io_s(FullAdder_189_io_s),
    .io_co(FullAdder_189_io_co)
  );
  FullAdder FullAdder_190 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_190_io_a),
    .io_b(FullAdder_190_io_b),
    .io_ci(FullAdder_190_io_ci),
    .io_s(FullAdder_190_io_s),
    .io_co(FullAdder_190_io_co)
  );
  FullAdder FullAdder_191 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_191_io_a),
    .io_b(FullAdder_191_io_b),
    .io_ci(FullAdder_191_io_ci),
    .io_s(FullAdder_191_io_s),
    .io_co(FullAdder_191_io_co)
  );
  FullAdder FullAdder_192 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_192_io_a),
    .io_b(FullAdder_192_io_b),
    .io_ci(FullAdder_192_io_ci),
    .io_s(FullAdder_192_io_s),
    .io_co(FullAdder_192_io_co)
  );
  FullAdder FullAdder_193 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_193_io_a),
    .io_b(FullAdder_193_io_b),
    .io_ci(FullAdder_193_io_ci),
    .io_s(FullAdder_193_io_s),
    .io_co(FullAdder_193_io_co)
  );
  FullAdder FullAdder_194 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_194_io_a),
    .io_b(FullAdder_194_io_b),
    .io_ci(FullAdder_194_io_ci),
    .io_s(FullAdder_194_io_s),
    .io_co(FullAdder_194_io_co)
  );
  FullAdder FullAdder_195 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_195_io_a),
    .io_b(FullAdder_195_io_b),
    .io_ci(FullAdder_195_io_ci),
    .io_s(FullAdder_195_io_s),
    .io_co(FullAdder_195_io_co)
  );
  FullAdder FullAdder_196 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_196_io_a),
    .io_b(FullAdder_196_io_b),
    .io_ci(FullAdder_196_io_ci),
    .io_s(FullAdder_196_io_s),
    .io_co(FullAdder_196_io_co)
  );
  FullAdder FullAdder_197 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_197_io_a),
    .io_b(FullAdder_197_io_b),
    .io_ci(FullAdder_197_io_ci),
    .io_s(FullAdder_197_io_s),
    .io_co(FullAdder_197_io_co)
  );
  FullAdder FullAdder_198 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_198_io_a),
    .io_b(FullAdder_198_io_b),
    .io_ci(FullAdder_198_io_ci),
    .io_s(FullAdder_198_io_s),
    .io_co(FullAdder_198_io_co)
  );
  FullAdder FullAdder_199 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_199_io_a),
    .io_b(FullAdder_199_io_b),
    .io_ci(FullAdder_199_io_ci),
    .io_s(FullAdder_199_io_s),
    .io_co(FullAdder_199_io_co)
  );
  FullAdder FullAdder_200 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_200_io_a),
    .io_b(FullAdder_200_io_b),
    .io_ci(FullAdder_200_io_ci),
    .io_s(FullAdder_200_io_s),
    .io_co(FullAdder_200_io_co)
  );
  HalfAdder HalfAdder_3 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_3_io_a),
    .io_b(HalfAdder_3_io_b),
    .io_s(HalfAdder_3_io_s),
    .io_co(HalfAdder_3_io_co)
  );
  HalfAdder HalfAdder_4 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_4_io_a),
    .io_b(HalfAdder_4_io_b),
    .io_s(HalfAdder_4_io_s),
    .io_co(HalfAdder_4_io_co)
  );
  HalfAdder HalfAdder_5 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_5_io_a),
    .io_b(HalfAdder_5_io_b),
    .io_s(HalfAdder_5_io_s),
    .io_co(HalfAdder_5_io_co)
  );
  FullAdder FullAdder_201 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_201_io_a),
    .io_b(FullAdder_201_io_b),
    .io_ci(FullAdder_201_io_ci),
    .io_s(FullAdder_201_io_s),
    .io_co(FullAdder_201_io_co)
  );
  FullAdder FullAdder_202 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_202_io_a),
    .io_b(FullAdder_202_io_b),
    .io_ci(FullAdder_202_io_ci),
    .io_s(FullAdder_202_io_s),
    .io_co(FullAdder_202_io_co)
  );
  FullAdder FullAdder_203 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_203_io_a),
    .io_b(FullAdder_203_io_b),
    .io_ci(FullAdder_203_io_ci),
    .io_s(FullAdder_203_io_s),
    .io_co(FullAdder_203_io_co)
  );
  FullAdder FullAdder_204 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_204_io_a),
    .io_b(FullAdder_204_io_b),
    .io_ci(FullAdder_204_io_ci),
    .io_s(FullAdder_204_io_s),
    .io_co(FullAdder_204_io_co)
  );
  FullAdder FullAdder_205 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_205_io_a),
    .io_b(FullAdder_205_io_b),
    .io_ci(FullAdder_205_io_ci),
    .io_s(FullAdder_205_io_s),
    .io_co(FullAdder_205_io_co)
  );
  FullAdder FullAdder_206 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_206_io_a),
    .io_b(FullAdder_206_io_b),
    .io_ci(FullAdder_206_io_ci),
    .io_s(FullAdder_206_io_s),
    .io_co(FullAdder_206_io_co)
  );
  FullAdder FullAdder_207 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_207_io_a),
    .io_b(FullAdder_207_io_b),
    .io_ci(FullAdder_207_io_ci),
    .io_s(FullAdder_207_io_s),
    .io_co(FullAdder_207_io_co)
  );
  FullAdder FullAdder_208 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_208_io_a),
    .io_b(FullAdder_208_io_b),
    .io_ci(FullAdder_208_io_ci),
    .io_s(FullAdder_208_io_s),
    .io_co(FullAdder_208_io_co)
  );
  FullAdder FullAdder_209 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_209_io_a),
    .io_b(FullAdder_209_io_b),
    .io_ci(FullAdder_209_io_ci),
    .io_s(FullAdder_209_io_s),
    .io_co(FullAdder_209_io_co)
  );
  FullAdder FullAdder_210 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_210_io_a),
    .io_b(FullAdder_210_io_b),
    .io_ci(FullAdder_210_io_ci),
    .io_s(FullAdder_210_io_s),
    .io_co(FullAdder_210_io_co)
  );
  FullAdder FullAdder_211 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_211_io_a),
    .io_b(FullAdder_211_io_b),
    .io_ci(FullAdder_211_io_ci),
    .io_s(FullAdder_211_io_s),
    .io_co(FullAdder_211_io_co)
  );
  FullAdder FullAdder_212 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_212_io_a),
    .io_b(FullAdder_212_io_b),
    .io_ci(FullAdder_212_io_ci),
    .io_s(FullAdder_212_io_s),
    .io_co(FullAdder_212_io_co)
  );
  FullAdder FullAdder_213 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_213_io_a),
    .io_b(FullAdder_213_io_b),
    .io_ci(FullAdder_213_io_ci),
    .io_s(FullAdder_213_io_s),
    .io_co(FullAdder_213_io_co)
  );
  FullAdder FullAdder_214 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_214_io_a),
    .io_b(FullAdder_214_io_b),
    .io_ci(FullAdder_214_io_ci),
    .io_s(FullAdder_214_io_s),
    .io_co(FullAdder_214_io_co)
  );
  FullAdder FullAdder_215 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_215_io_a),
    .io_b(FullAdder_215_io_b),
    .io_ci(FullAdder_215_io_ci),
    .io_s(FullAdder_215_io_s),
    .io_co(FullAdder_215_io_co)
  );
  FullAdder FullAdder_216 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_216_io_a),
    .io_b(FullAdder_216_io_b),
    .io_ci(FullAdder_216_io_ci),
    .io_s(FullAdder_216_io_s),
    .io_co(FullAdder_216_io_co)
  );
  FullAdder FullAdder_217 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_217_io_a),
    .io_b(FullAdder_217_io_b),
    .io_ci(FullAdder_217_io_ci),
    .io_s(FullAdder_217_io_s),
    .io_co(FullAdder_217_io_co)
  );
  FullAdder FullAdder_218 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_218_io_a),
    .io_b(FullAdder_218_io_b),
    .io_ci(FullAdder_218_io_ci),
    .io_s(FullAdder_218_io_s),
    .io_co(FullAdder_218_io_co)
  );
  FullAdder FullAdder_219 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_219_io_a),
    .io_b(FullAdder_219_io_b),
    .io_ci(FullAdder_219_io_ci),
    .io_s(FullAdder_219_io_s),
    .io_co(FullAdder_219_io_co)
  );
  FullAdder FullAdder_220 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_220_io_a),
    .io_b(FullAdder_220_io_b),
    .io_ci(FullAdder_220_io_ci),
    .io_s(FullAdder_220_io_s),
    .io_co(FullAdder_220_io_co)
  );
  FullAdder FullAdder_221 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_221_io_a),
    .io_b(FullAdder_221_io_b),
    .io_ci(FullAdder_221_io_ci),
    .io_s(FullAdder_221_io_s),
    .io_co(FullAdder_221_io_co)
  );
  FullAdder FullAdder_222 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_222_io_a),
    .io_b(FullAdder_222_io_b),
    .io_ci(FullAdder_222_io_ci),
    .io_s(FullAdder_222_io_s),
    .io_co(FullAdder_222_io_co)
  );
  FullAdder FullAdder_223 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_223_io_a),
    .io_b(FullAdder_223_io_b),
    .io_ci(FullAdder_223_io_ci),
    .io_s(FullAdder_223_io_s),
    .io_co(FullAdder_223_io_co)
  );
  FullAdder FullAdder_224 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_224_io_a),
    .io_b(FullAdder_224_io_b),
    .io_ci(FullAdder_224_io_ci),
    .io_s(FullAdder_224_io_s),
    .io_co(FullAdder_224_io_co)
  );
  FullAdder FullAdder_225 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_225_io_a),
    .io_b(FullAdder_225_io_b),
    .io_ci(FullAdder_225_io_ci),
    .io_s(FullAdder_225_io_s),
    .io_co(FullAdder_225_io_co)
  );
  FullAdder FullAdder_226 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_226_io_a),
    .io_b(FullAdder_226_io_b),
    .io_ci(FullAdder_226_io_ci),
    .io_s(FullAdder_226_io_s),
    .io_co(FullAdder_226_io_co)
  );
  FullAdder FullAdder_227 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_227_io_a),
    .io_b(FullAdder_227_io_b),
    .io_ci(FullAdder_227_io_ci),
    .io_s(FullAdder_227_io_s),
    .io_co(FullAdder_227_io_co)
  );
  FullAdder FullAdder_228 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_228_io_a),
    .io_b(FullAdder_228_io_b),
    .io_ci(FullAdder_228_io_ci),
    .io_s(FullAdder_228_io_s),
    .io_co(FullAdder_228_io_co)
  );
  FullAdder FullAdder_229 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_229_io_a),
    .io_b(FullAdder_229_io_b),
    .io_ci(FullAdder_229_io_ci),
    .io_s(FullAdder_229_io_s),
    .io_co(FullAdder_229_io_co)
  );
  FullAdder FullAdder_230 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_230_io_a),
    .io_b(FullAdder_230_io_b),
    .io_ci(FullAdder_230_io_ci),
    .io_s(FullAdder_230_io_s),
    .io_co(FullAdder_230_io_co)
  );
  FullAdder FullAdder_231 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_231_io_a),
    .io_b(FullAdder_231_io_b),
    .io_ci(FullAdder_231_io_ci),
    .io_s(FullAdder_231_io_s),
    .io_co(FullAdder_231_io_co)
  );
  FullAdder FullAdder_232 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_232_io_a),
    .io_b(FullAdder_232_io_b),
    .io_ci(FullAdder_232_io_ci),
    .io_s(FullAdder_232_io_s),
    .io_co(FullAdder_232_io_co)
  );
  FullAdder FullAdder_233 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_233_io_a),
    .io_b(FullAdder_233_io_b),
    .io_ci(FullAdder_233_io_ci),
    .io_s(FullAdder_233_io_s),
    .io_co(FullAdder_233_io_co)
  );
  FullAdder FullAdder_234 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_234_io_a),
    .io_b(FullAdder_234_io_b),
    .io_ci(FullAdder_234_io_ci),
    .io_s(FullAdder_234_io_s),
    .io_co(FullAdder_234_io_co)
  );
  FullAdder FullAdder_235 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_235_io_a),
    .io_b(FullAdder_235_io_b),
    .io_ci(FullAdder_235_io_ci),
    .io_s(FullAdder_235_io_s),
    .io_co(FullAdder_235_io_co)
  );
  FullAdder FullAdder_236 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_236_io_a),
    .io_b(FullAdder_236_io_b),
    .io_ci(FullAdder_236_io_ci),
    .io_s(FullAdder_236_io_s),
    .io_co(FullAdder_236_io_co)
  );
  FullAdder FullAdder_237 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_237_io_a),
    .io_b(FullAdder_237_io_b),
    .io_ci(FullAdder_237_io_ci),
    .io_s(FullAdder_237_io_s),
    .io_co(FullAdder_237_io_co)
  );
  FullAdder FullAdder_238 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_238_io_a),
    .io_b(FullAdder_238_io_b),
    .io_ci(FullAdder_238_io_ci),
    .io_s(FullAdder_238_io_s),
    .io_co(FullAdder_238_io_co)
  );
  FullAdder FullAdder_239 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_239_io_a),
    .io_b(FullAdder_239_io_b),
    .io_ci(FullAdder_239_io_ci),
    .io_s(FullAdder_239_io_s),
    .io_co(FullAdder_239_io_co)
  );
  FullAdder FullAdder_240 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_240_io_a),
    .io_b(FullAdder_240_io_b),
    .io_ci(FullAdder_240_io_ci),
    .io_s(FullAdder_240_io_s),
    .io_co(FullAdder_240_io_co)
  );
  FullAdder FullAdder_241 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_241_io_a),
    .io_b(FullAdder_241_io_b),
    .io_ci(FullAdder_241_io_ci),
    .io_s(FullAdder_241_io_s),
    .io_co(FullAdder_241_io_co)
  );
  FullAdder FullAdder_242 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_242_io_a),
    .io_b(FullAdder_242_io_b),
    .io_ci(FullAdder_242_io_ci),
    .io_s(FullAdder_242_io_s),
    .io_co(FullAdder_242_io_co)
  );
  FullAdder FullAdder_243 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_243_io_a),
    .io_b(FullAdder_243_io_b),
    .io_ci(FullAdder_243_io_ci),
    .io_s(FullAdder_243_io_s),
    .io_co(FullAdder_243_io_co)
  );
  FullAdder FullAdder_244 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_244_io_a),
    .io_b(FullAdder_244_io_b),
    .io_ci(FullAdder_244_io_ci),
    .io_s(FullAdder_244_io_s),
    .io_co(FullAdder_244_io_co)
  );
  FullAdder FullAdder_245 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_245_io_a),
    .io_b(FullAdder_245_io_b),
    .io_ci(FullAdder_245_io_ci),
    .io_s(FullAdder_245_io_s),
    .io_co(FullAdder_245_io_co)
  );
  FullAdder FullAdder_246 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_246_io_a),
    .io_b(FullAdder_246_io_b),
    .io_ci(FullAdder_246_io_ci),
    .io_s(FullAdder_246_io_s),
    .io_co(FullAdder_246_io_co)
  );
  FullAdder FullAdder_247 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_247_io_a),
    .io_b(FullAdder_247_io_b),
    .io_ci(FullAdder_247_io_ci),
    .io_s(FullAdder_247_io_s),
    .io_co(FullAdder_247_io_co)
  );
  FullAdder FullAdder_248 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_248_io_a),
    .io_b(FullAdder_248_io_b),
    .io_ci(FullAdder_248_io_ci),
    .io_s(FullAdder_248_io_s),
    .io_co(FullAdder_248_io_co)
  );
  FullAdder FullAdder_249 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_249_io_a),
    .io_b(FullAdder_249_io_b),
    .io_ci(FullAdder_249_io_ci),
    .io_s(FullAdder_249_io_s),
    .io_co(FullAdder_249_io_co)
  );
  FullAdder FullAdder_250 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_250_io_a),
    .io_b(FullAdder_250_io_b),
    .io_ci(FullAdder_250_io_ci),
    .io_s(FullAdder_250_io_s),
    .io_co(FullAdder_250_io_co)
  );
  FullAdder FullAdder_251 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_251_io_a),
    .io_b(FullAdder_251_io_b),
    .io_ci(FullAdder_251_io_ci),
    .io_s(FullAdder_251_io_s),
    .io_co(FullAdder_251_io_co)
  );
  FullAdder FullAdder_252 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_252_io_a),
    .io_b(FullAdder_252_io_b),
    .io_ci(FullAdder_252_io_ci),
    .io_s(FullAdder_252_io_s),
    .io_co(FullAdder_252_io_co)
  );
  FullAdder FullAdder_253 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_253_io_a),
    .io_b(FullAdder_253_io_b),
    .io_ci(FullAdder_253_io_ci),
    .io_s(FullAdder_253_io_s),
    .io_co(FullAdder_253_io_co)
  );
  FullAdder FullAdder_254 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_254_io_a),
    .io_b(FullAdder_254_io_b),
    .io_ci(FullAdder_254_io_ci),
    .io_s(FullAdder_254_io_s),
    .io_co(FullAdder_254_io_co)
  );
  FullAdder FullAdder_255 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_255_io_a),
    .io_b(FullAdder_255_io_b),
    .io_ci(FullAdder_255_io_ci),
    .io_s(FullAdder_255_io_s),
    .io_co(FullAdder_255_io_co)
  );
  FullAdder FullAdder_256 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_256_io_a),
    .io_b(FullAdder_256_io_b),
    .io_ci(FullAdder_256_io_ci),
    .io_s(FullAdder_256_io_s),
    .io_co(FullAdder_256_io_co)
  );
  FullAdder FullAdder_257 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_257_io_a),
    .io_b(FullAdder_257_io_b),
    .io_ci(FullAdder_257_io_ci),
    .io_s(FullAdder_257_io_s),
    .io_co(FullAdder_257_io_co)
  );
  FullAdder FullAdder_258 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_258_io_a),
    .io_b(FullAdder_258_io_b),
    .io_ci(FullAdder_258_io_ci),
    .io_s(FullAdder_258_io_s),
    .io_co(FullAdder_258_io_co)
  );
  FullAdder FullAdder_259 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_259_io_a),
    .io_b(FullAdder_259_io_b),
    .io_ci(FullAdder_259_io_ci),
    .io_s(FullAdder_259_io_s),
    .io_co(FullAdder_259_io_co)
  );
  FullAdder FullAdder_260 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_260_io_a),
    .io_b(FullAdder_260_io_b),
    .io_ci(FullAdder_260_io_ci),
    .io_s(FullAdder_260_io_s),
    .io_co(FullAdder_260_io_co)
  );
  FullAdder FullAdder_261 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_261_io_a),
    .io_b(FullAdder_261_io_b),
    .io_ci(FullAdder_261_io_ci),
    .io_s(FullAdder_261_io_s),
    .io_co(FullAdder_261_io_co)
  );
  FullAdder FullAdder_262 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_262_io_a),
    .io_b(FullAdder_262_io_b),
    .io_ci(FullAdder_262_io_ci),
    .io_s(FullAdder_262_io_s),
    .io_co(FullAdder_262_io_co)
  );
  FullAdder FullAdder_263 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_263_io_a),
    .io_b(FullAdder_263_io_b),
    .io_ci(FullAdder_263_io_ci),
    .io_s(FullAdder_263_io_s),
    .io_co(FullAdder_263_io_co)
  );
  FullAdder FullAdder_264 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_264_io_a),
    .io_b(FullAdder_264_io_b),
    .io_ci(FullAdder_264_io_ci),
    .io_s(FullAdder_264_io_s),
    .io_co(FullAdder_264_io_co)
  );
  FullAdder FullAdder_265 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_265_io_a),
    .io_b(FullAdder_265_io_b),
    .io_ci(FullAdder_265_io_ci),
    .io_s(FullAdder_265_io_s),
    .io_co(FullAdder_265_io_co)
  );
  FullAdder FullAdder_266 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_266_io_a),
    .io_b(FullAdder_266_io_b),
    .io_ci(FullAdder_266_io_ci),
    .io_s(FullAdder_266_io_s),
    .io_co(FullAdder_266_io_co)
  );
  FullAdder FullAdder_267 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_267_io_a),
    .io_b(FullAdder_267_io_b),
    .io_ci(FullAdder_267_io_ci),
    .io_s(FullAdder_267_io_s),
    .io_co(FullAdder_267_io_co)
  );
  FullAdder FullAdder_268 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_268_io_a),
    .io_b(FullAdder_268_io_b),
    .io_ci(FullAdder_268_io_ci),
    .io_s(FullAdder_268_io_s),
    .io_co(FullAdder_268_io_co)
  );
  FullAdder FullAdder_269 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_269_io_a),
    .io_b(FullAdder_269_io_b),
    .io_ci(FullAdder_269_io_ci),
    .io_s(FullAdder_269_io_s),
    .io_co(FullAdder_269_io_co)
  );
  FullAdder FullAdder_270 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_270_io_a),
    .io_b(FullAdder_270_io_b),
    .io_ci(FullAdder_270_io_ci),
    .io_s(FullAdder_270_io_s),
    .io_co(FullAdder_270_io_co)
  );
  FullAdder FullAdder_271 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_271_io_a),
    .io_b(FullAdder_271_io_b),
    .io_ci(FullAdder_271_io_ci),
    .io_s(FullAdder_271_io_s),
    .io_co(FullAdder_271_io_co)
  );
  FullAdder FullAdder_272 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_272_io_a),
    .io_b(FullAdder_272_io_b),
    .io_ci(FullAdder_272_io_ci),
    .io_s(FullAdder_272_io_s),
    .io_co(FullAdder_272_io_co)
  );
  FullAdder FullAdder_273 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_273_io_a),
    .io_b(FullAdder_273_io_b),
    .io_ci(FullAdder_273_io_ci),
    .io_s(FullAdder_273_io_s),
    .io_co(FullAdder_273_io_co)
  );
  FullAdder FullAdder_274 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_274_io_a),
    .io_b(FullAdder_274_io_b),
    .io_ci(FullAdder_274_io_ci),
    .io_s(FullAdder_274_io_s),
    .io_co(FullAdder_274_io_co)
  );
  FullAdder FullAdder_275 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_275_io_a),
    .io_b(FullAdder_275_io_b),
    .io_ci(FullAdder_275_io_ci),
    .io_s(FullAdder_275_io_s),
    .io_co(FullAdder_275_io_co)
  );
  FullAdder FullAdder_276 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_276_io_a),
    .io_b(FullAdder_276_io_b),
    .io_ci(FullAdder_276_io_ci),
    .io_s(FullAdder_276_io_s),
    .io_co(FullAdder_276_io_co)
  );
  FullAdder FullAdder_277 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_277_io_a),
    .io_b(FullAdder_277_io_b),
    .io_ci(FullAdder_277_io_ci),
    .io_s(FullAdder_277_io_s),
    .io_co(FullAdder_277_io_co)
  );
  FullAdder FullAdder_278 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_278_io_a),
    .io_b(FullAdder_278_io_b),
    .io_ci(FullAdder_278_io_ci),
    .io_s(FullAdder_278_io_s),
    .io_co(FullAdder_278_io_co)
  );
  FullAdder FullAdder_279 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_279_io_a),
    .io_b(FullAdder_279_io_b),
    .io_ci(FullAdder_279_io_ci),
    .io_s(FullAdder_279_io_s),
    .io_co(FullAdder_279_io_co)
  );
  FullAdder FullAdder_280 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_280_io_a),
    .io_b(FullAdder_280_io_b),
    .io_ci(FullAdder_280_io_ci),
    .io_s(FullAdder_280_io_s),
    .io_co(FullAdder_280_io_co)
  );
  FullAdder FullAdder_281 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_281_io_a),
    .io_b(FullAdder_281_io_b),
    .io_ci(FullAdder_281_io_ci),
    .io_s(FullAdder_281_io_s),
    .io_co(FullAdder_281_io_co)
  );
  FullAdder FullAdder_282 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_282_io_a),
    .io_b(FullAdder_282_io_b),
    .io_ci(FullAdder_282_io_ci),
    .io_s(FullAdder_282_io_s),
    .io_co(FullAdder_282_io_co)
  );
  FullAdder FullAdder_283 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_283_io_a),
    .io_b(FullAdder_283_io_b),
    .io_ci(FullAdder_283_io_ci),
    .io_s(FullAdder_283_io_s),
    .io_co(FullAdder_283_io_co)
  );
  FullAdder FullAdder_284 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_284_io_a),
    .io_b(FullAdder_284_io_b),
    .io_ci(FullAdder_284_io_ci),
    .io_s(FullAdder_284_io_s),
    .io_co(FullAdder_284_io_co)
  );
  FullAdder FullAdder_285 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_285_io_a),
    .io_b(FullAdder_285_io_b),
    .io_ci(FullAdder_285_io_ci),
    .io_s(FullAdder_285_io_s),
    .io_co(FullAdder_285_io_co)
  );
  FullAdder FullAdder_286 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_286_io_a),
    .io_b(FullAdder_286_io_b),
    .io_ci(FullAdder_286_io_ci),
    .io_s(FullAdder_286_io_s),
    .io_co(FullAdder_286_io_co)
  );
  FullAdder FullAdder_287 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_287_io_a),
    .io_b(FullAdder_287_io_b),
    .io_ci(FullAdder_287_io_ci),
    .io_s(FullAdder_287_io_s),
    .io_co(FullAdder_287_io_co)
  );
  FullAdder FullAdder_288 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_288_io_a),
    .io_b(FullAdder_288_io_b),
    .io_ci(FullAdder_288_io_ci),
    .io_s(FullAdder_288_io_s),
    .io_co(FullAdder_288_io_co)
  );
  FullAdder FullAdder_289 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_289_io_a),
    .io_b(FullAdder_289_io_b),
    .io_ci(FullAdder_289_io_ci),
    .io_s(FullAdder_289_io_s),
    .io_co(FullAdder_289_io_co)
  );
  FullAdder FullAdder_290 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_290_io_a),
    .io_b(FullAdder_290_io_b),
    .io_ci(FullAdder_290_io_ci),
    .io_s(FullAdder_290_io_s),
    .io_co(FullAdder_290_io_co)
  );
  FullAdder FullAdder_291 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_291_io_a),
    .io_b(FullAdder_291_io_b),
    .io_ci(FullAdder_291_io_ci),
    .io_s(FullAdder_291_io_s),
    .io_co(FullAdder_291_io_co)
  );
  FullAdder FullAdder_292 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_292_io_a),
    .io_b(FullAdder_292_io_b),
    .io_ci(FullAdder_292_io_ci),
    .io_s(FullAdder_292_io_s),
    .io_co(FullAdder_292_io_co)
  );
  FullAdder FullAdder_293 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_293_io_a),
    .io_b(FullAdder_293_io_b),
    .io_ci(FullAdder_293_io_ci),
    .io_s(FullAdder_293_io_s),
    .io_co(FullAdder_293_io_co)
  );
  FullAdder FullAdder_294 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_294_io_a),
    .io_b(FullAdder_294_io_b),
    .io_ci(FullAdder_294_io_ci),
    .io_s(FullAdder_294_io_s),
    .io_co(FullAdder_294_io_co)
  );
  FullAdder FullAdder_295 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_295_io_a),
    .io_b(FullAdder_295_io_b),
    .io_ci(FullAdder_295_io_ci),
    .io_s(FullAdder_295_io_s),
    .io_co(FullAdder_295_io_co)
  );
  FullAdder FullAdder_296 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_296_io_a),
    .io_b(FullAdder_296_io_b),
    .io_ci(FullAdder_296_io_ci),
    .io_s(FullAdder_296_io_s),
    .io_co(FullAdder_296_io_co)
  );
  FullAdder FullAdder_297 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_297_io_a),
    .io_b(FullAdder_297_io_b),
    .io_ci(FullAdder_297_io_ci),
    .io_s(FullAdder_297_io_s),
    .io_co(FullAdder_297_io_co)
  );
  FullAdder FullAdder_298 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_298_io_a),
    .io_b(FullAdder_298_io_b),
    .io_ci(FullAdder_298_io_ci),
    .io_s(FullAdder_298_io_s),
    .io_co(FullAdder_298_io_co)
  );
  FullAdder FullAdder_299 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_299_io_a),
    .io_b(FullAdder_299_io_b),
    .io_ci(FullAdder_299_io_ci),
    .io_s(FullAdder_299_io_s),
    .io_co(FullAdder_299_io_co)
  );
  FullAdder FullAdder_300 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_300_io_a),
    .io_b(FullAdder_300_io_b),
    .io_ci(FullAdder_300_io_ci),
    .io_s(FullAdder_300_io_s),
    .io_co(FullAdder_300_io_co)
  );
  FullAdder FullAdder_301 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_301_io_a),
    .io_b(FullAdder_301_io_b),
    .io_ci(FullAdder_301_io_ci),
    .io_s(FullAdder_301_io_s),
    .io_co(FullAdder_301_io_co)
  );
  FullAdder FullAdder_302 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_302_io_a),
    .io_b(FullAdder_302_io_b),
    .io_ci(FullAdder_302_io_ci),
    .io_s(FullAdder_302_io_s),
    .io_co(FullAdder_302_io_co)
  );
  FullAdder FullAdder_303 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_303_io_a),
    .io_b(FullAdder_303_io_b),
    .io_ci(FullAdder_303_io_ci),
    .io_s(FullAdder_303_io_s),
    .io_co(FullAdder_303_io_co)
  );
  FullAdder FullAdder_304 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_304_io_a),
    .io_b(FullAdder_304_io_b),
    .io_ci(FullAdder_304_io_ci),
    .io_s(FullAdder_304_io_s),
    .io_co(FullAdder_304_io_co)
  );
  FullAdder FullAdder_305 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_305_io_a),
    .io_b(FullAdder_305_io_b),
    .io_ci(FullAdder_305_io_ci),
    .io_s(FullAdder_305_io_s),
    .io_co(FullAdder_305_io_co)
  );
  FullAdder FullAdder_306 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_306_io_a),
    .io_b(FullAdder_306_io_b),
    .io_ci(FullAdder_306_io_ci),
    .io_s(FullAdder_306_io_s),
    .io_co(FullAdder_306_io_co)
  );
  FullAdder FullAdder_307 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_307_io_a),
    .io_b(FullAdder_307_io_b),
    .io_ci(FullAdder_307_io_ci),
    .io_s(FullAdder_307_io_s),
    .io_co(FullAdder_307_io_co)
  );
  FullAdder FullAdder_308 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_308_io_a),
    .io_b(FullAdder_308_io_b),
    .io_ci(FullAdder_308_io_ci),
    .io_s(FullAdder_308_io_s),
    .io_co(FullAdder_308_io_co)
  );
  FullAdder FullAdder_309 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_309_io_a),
    .io_b(FullAdder_309_io_b),
    .io_ci(FullAdder_309_io_ci),
    .io_s(FullAdder_309_io_s),
    .io_co(FullAdder_309_io_co)
  );
  FullAdder FullAdder_310 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_310_io_a),
    .io_b(FullAdder_310_io_b),
    .io_ci(FullAdder_310_io_ci),
    .io_s(FullAdder_310_io_s),
    .io_co(FullAdder_310_io_co)
  );
  FullAdder FullAdder_311 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_311_io_a),
    .io_b(FullAdder_311_io_b),
    .io_ci(FullAdder_311_io_ci),
    .io_s(FullAdder_311_io_s),
    .io_co(FullAdder_311_io_co)
  );
  FullAdder FullAdder_312 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_312_io_a),
    .io_b(FullAdder_312_io_b),
    .io_ci(FullAdder_312_io_ci),
    .io_s(FullAdder_312_io_s),
    .io_co(FullAdder_312_io_co)
  );
  FullAdder FullAdder_313 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_313_io_a),
    .io_b(FullAdder_313_io_b),
    .io_ci(FullAdder_313_io_ci),
    .io_s(FullAdder_313_io_s),
    .io_co(FullAdder_313_io_co)
  );
  FullAdder FullAdder_314 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_314_io_a),
    .io_b(FullAdder_314_io_b),
    .io_ci(FullAdder_314_io_ci),
    .io_s(FullAdder_314_io_s),
    .io_co(FullAdder_314_io_co)
  );
  FullAdder FullAdder_315 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_315_io_a),
    .io_b(FullAdder_315_io_b),
    .io_ci(FullAdder_315_io_ci),
    .io_s(FullAdder_315_io_s),
    .io_co(FullAdder_315_io_co)
  );
  FullAdder FullAdder_316 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_316_io_a),
    .io_b(FullAdder_316_io_b),
    .io_ci(FullAdder_316_io_ci),
    .io_s(FullAdder_316_io_s),
    .io_co(FullAdder_316_io_co)
  );
  FullAdder FullAdder_317 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_317_io_a),
    .io_b(FullAdder_317_io_b),
    .io_ci(FullAdder_317_io_ci),
    .io_s(FullAdder_317_io_s),
    .io_co(FullAdder_317_io_co)
  );
  FullAdder FullAdder_318 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_318_io_a),
    .io_b(FullAdder_318_io_b),
    .io_ci(FullAdder_318_io_ci),
    .io_s(FullAdder_318_io_s),
    .io_co(FullAdder_318_io_co)
  );
  FullAdder FullAdder_319 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_319_io_a),
    .io_b(FullAdder_319_io_b),
    .io_ci(FullAdder_319_io_ci),
    .io_s(FullAdder_319_io_s),
    .io_co(FullAdder_319_io_co)
  );
  FullAdder FullAdder_320 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_320_io_a),
    .io_b(FullAdder_320_io_b),
    .io_ci(FullAdder_320_io_ci),
    .io_s(FullAdder_320_io_s),
    .io_co(FullAdder_320_io_co)
  );
  FullAdder FullAdder_321 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_321_io_a),
    .io_b(FullAdder_321_io_b),
    .io_ci(FullAdder_321_io_ci),
    .io_s(FullAdder_321_io_s),
    .io_co(FullAdder_321_io_co)
  );
  FullAdder FullAdder_322 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_322_io_a),
    .io_b(FullAdder_322_io_b),
    .io_ci(FullAdder_322_io_ci),
    .io_s(FullAdder_322_io_s),
    .io_co(FullAdder_322_io_co)
  );
  FullAdder FullAdder_323 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_323_io_a),
    .io_b(FullAdder_323_io_b),
    .io_ci(FullAdder_323_io_ci),
    .io_s(FullAdder_323_io_s),
    .io_co(FullAdder_323_io_co)
  );
  FullAdder FullAdder_324 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_324_io_a),
    .io_b(FullAdder_324_io_b),
    .io_ci(FullAdder_324_io_ci),
    .io_s(FullAdder_324_io_s),
    .io_co(FullAdder_324_io_co)
  );
  FullAdder FullAdder_325 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_325_io_a),
    .io_b(FullAdder_325_io_b),
    .io_ci(FullAdder_325_io_ci),
    .io_s(FullAdder_325_io_s),
    .io_co(FullAdder_325_io_co)
  );
  FullAdder FullAdder_326 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_326_io_a),
    .io_b(FullAdder_326_io_b),
    .io_ci(FullAdder_326_io_ci),
    .io_s(FullAdder_326_io_s),
    .io_co(FullAdder_326_io_co)
  );
  FullAdder FullAdder_327 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_327_io_a),
    .io_b(FullAdder_327_io_b),
    .io_ci(FullAdder_327_io_ci),
    .io_s(FullAdder_327_io_s),
    .io_co(FullAdder_327_io_co)
  );
  FullAdder FullAdder_328 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_328_io_a),
    .io_b(FullAdder_328_io_b),
    .io_ci(FullAdder_328_io_ci),
    .io_s(FullAdder_328_io_s),
    .io_co(FullAdder_328_io_co)
  );
  FullAdder FullAdder_329 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_329_io_a),
    .io_b(FullAdder_329_io_b),
    .io_ci(FullAdder_329_io_ci),
    .io_s(FullAdder_329_io_s),
    .io_co(FullAdder_329_io_co)
  );
  FullAdder FullAdder_330 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_330_io_a),
    .io_b(FullAdder_330_io_b),
    .io_ci(FullAdder_330_io_ci),
    .io_s(FullAdder_330_io_s),
    .io_co(FullAdder_330_io_co)
  );
  FullAdder FullAdder_331 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_331_io_a),
    .io_b(FullAdder_331_io_b),
    .io_ci(FullAdder_331_io_ci),
    .io_s(FullAdder_331_io_s),
    .io_co(FullAdder_331_io_co)
  );
  FullAdder FullAdder_332 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_332_io_a),
    .io_b(FullAdder_332_io_b),
    .io_ci(FullAdder_332_io_ci),
    .io_s(FullAdder_332_io_s),
    .io_co(FullAdder_332_io_co)
  );
  FullAdder FullAdder_333 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_333_io_a),
    .io_b(FullAdder_333_io_b),
    .io_ci(FullAdder_333_io_ci),
    .io_s(FullAdder_333_io_s),
    .io_co(FullAdder_333_io_co)
  );
  FullAdder FullAdder_334 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_334_io_a),
    .io_b(FullAdder_334_io_b),
    .io_ci(FullAdder_334_io_ci),
    .io_s(FullAdder_334_io_s),
    .io_co(FullAdder_334_io_co)
  );
  FullAdder FullAdder_335 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_335_io_a),
    .io_b(FullAdder_335_io_b),
    .io_ci(FullAdder_335_io_ci),
    .io_s(FullAdder_335_io_s),
    .io_co(FullAdder_335_io_co)
  );
  FullAdder FullAdder_336 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_336_io_a),
    .io_b(FullAdder_336_io_b),
    .io_ci(FullAdder_336_io_ci),
    .io_s(FullAdder_336_io_s),
    .io_co(FullAdder_336_io_co)
  );
  FullAdder FullAdder_337 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_337_io_a),
    .io_b(FullAdder_337_io_b),
    .io_ci(FullAdder_337_io_ci),
    .io_s(FullAdder_337_io_s),
    .io_co(FullAdder_337_io_co)
  );
  FullAdder FullAdder_338 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_338_io_a),
    .io_b(FullAdder_338_io_b),
    .io_ci(FullAdder_338_io_ci),
    .io_s(FullAdder_338_io_s),
    .io_co(FullAdder_338_io_co)
  );
  FullAdder FullAdder_339 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_339_io_a),
    .io_b(FullAdder_339_io_b),
    .io_ci(FullAdder_339_io_ci),
    .io_s(FullAdder_339_io_s),
    .io_co(FullAdder_339_io_co)
  );
  FullAdder FullAdder_340 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_340_io_a),
    .io_b(FullAdder_340_io_b),
    .io_ci(FullAdder_340_io_ci),
    .io_s(FullAdder_340_io_s),
    .io_co(FullAdder_340_io_co)
  );
  FullAdder FullAdder_341 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_341_io_a),
    .io_b(FullAdder_341_io_b),
    .io_ci(FullAdder_341_io_ci),
    .io_s(FullAdder_341_io_s),
    .io_co(FullAdder_341_io_co)
  );
  FullAdder FullAdder_342 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_342_io_a),
    .io_b(FullAdder_342_io_b),
    .io_ci(FullAdder_342_io_ci),
    .io_s(FullAdder_342_io_s),
    .io_co(FullAdder_342_io_co)
  );
  FullAdder FullAdder_343 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_343_io_a),
    .io_b(FullAdder_343_io_b),
    .io_ci(FullAdder_343_io_ci),
    .io_s(FullAdder_343_io_s),
    .io_co(FullAdder_343_io_co)
  );
  FullAdder FullAdder_344 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_344_io_a),
    .io_b(FullAdder_344_io_b),
    .io_ci(FullAdder_344_io_ci),
    .io_s(FullAdder_344_io_s),
    .io_co(FullAdder_344_io_co)
  );
  FullAdder FullAdder_345 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_345_io_a),
    .io_b(FullAdder_345_io_b),
    .io_ci(FullAdder_345_io_ci),
    .io_s(FullAdder_345_io_s),
    .io_co(FullAdder_345_io_co)
  );
  FullAdder FullAdder_346 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_346_io_a),
    .io_b(FullAdder_346_io_b),
    .io_ci(FullAdder_346_io_ci),
    .io_s(FullAdder_346_io_s),
    .io_co(FullAdder_346_io_co)
  );
  FullAdder FullAdder_347 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_347_io_a),
    .io_b(FullAdder_347_io_b),
    .io_ci(FullAdder_347_io_ci),
    .io_s(FullAdder_347_io_s),
    .io_co(FullAdder_347_io_co)
  );
  FullAdder FullAdder_348 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_348_io_a),
    .io_b(FullAdder_348_io_b),
    .io_ci(FullAdder_348_io_ci),
    .io_s(FullAdder_348_io_s),
    .io_co(FullAdder_348_io_co)
  );
  FullAdder FullAdder_349 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_349_io_a),
    .io_b(FullAdder_349_io_b),
    .io_ci(FullAdder_349_io_ci),
    .io_s(FullAdder_349_io_s),
    .io_co(FullAdder_349_io_co)
  );
  FullAdder FullAdder_350 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_350_io_a),
    .io_b(FullAdder_350_io_b),
    .io_ci(FullAdder_350_io_ci),
    .io_s(FullAdder_350_io_s),
    .io_co(FullAdder_350_io_co)
  );
  FullAdder FullAdder_351 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_351_io_a),
    .io_b(FullAdder_351_io_b),
    .io_ci(FullAdder_351_io_ci),
    .io_s(FullAdder_351_io_s),
    .io_co(FullAdder_351_io_co)
  );
  FullAdder FullAdder_352 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_352_io_a),
    .io_b(FullAdder_352_io_b),
    .io_ci(FullAdder_352_io_ci),
    .io_s(FullAdder_352_io_s),
    .io_co(FullAdder_352_io_co)
  );
  FullAdder FullAdder_353 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_353_io_a),
    .io_b(FullAdder_353_io_b),
    .io_ci(FullAdder_353_io_ci),
    .io_s(FullAdder_353_io_s),
    .io_co(FullAdder_353_io_co)
  );
  FullAdder FullAdder_354 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_354_io_a),
    .io_b(FullAdder_354_io_b),
    .io_ci(FullAdder_354_io_ci),
    .io_s(FullAdder_354_io_s),
    .io_co(FullAdder_354_io_co)
  );
  FullAdder FullAdder_355 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_355_io_a),
    .io_b(FullAdder_355_io_b),
    .io_ci(FullAdder_355_io_ci),
    .io_s(FullAdder_355_io_s),
    .io_co(FullAdder_355_io_co)
  );
  FullAdder FullAdder_356 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_356_io_a),
    .io_b(FullAdder_356_io_b),
    .io_ci(FullAdder_356_io_ci),
    .io_s(FullAdder_356_io_s),
    .io_co(FullAdder_356_io_co)
  );
  FullAdder FullAdder_357 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_357_io_a),
    .io_b(FullAdder_357_io_b),
    .io_ci(FullAdder_357_io_ci),
    .io_s(FullAdder_357_io_s),
    .io_co(FullAdder_357_io_co)
  );
  HalfAdder HalfAdder_6 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_6_io_a),
    .io_b(HalfAdder_6_io_b),
    .io_s(HalfAdder_6_io_s),
    .io_co(HalfAdder_6_io_co)
  );
  FullAdder FullAdder_358 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_358_io_a),
    .io_b(FullAdder_358_io_b),
    .io_ci(FullAdder_358_io_ci),
    .io_s(FullAdder_358_io_s),
    .io_co(FullAdder_358_io_co)
  );
  FullAdder FullAdder_359 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_359_io_a),
    .io_b(FullAdder_359_io_b),
    .io_ci(FullAdder_359_io_ci),
    .io_s(FullAdder_359_io_s),
    .io_co(FullAdder_359_io_co)
  );
  FullAdder FullAdder_360 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_360_io_a),
    .io_b(FullAdder_360_io_b),
    .io_ci(FullAdder_360_io_ci),
    .io_s(FullAdder_360_io_s),
    .io_co(FullAdder_360_io_co)
  );
  FullAdder FullAdder_361 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_361_io_a),
    .io_b(FullAdder_361_io_b),
    .io_ci(FullAdder_361_io_ci),
    .io_s(FullAdder_361_io_s),
    .io_co(FullAdder_361_io_co)
  );
  FullAdder FullAdder_362 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_362_io_a),
    .io_b(FullAdder_362_io_b),
    .io_ci(FullAdder_362_io_ci),
    .io_s(FullAdder_362_io_s),
    .io_co(FullAdder_362_io_co)
  );
  FullAdder FullAdder_363 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_363_io_a),
    .io_b(FullAdder_363_io_b),
    .io_ci(FullAdder_363_io_ci),
    .io_s(FullAdder_363_io_s),
    .io_co(FullAdder_363_io_co)
  );
  FullAdder FullAdder_364 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_364_io_a),
    .io_b(FullAdder_364_io_b),
    .io_ci(FullAdder_364_io_ci),
    .io_s(FullAdder_364_io_s),
    .io_co(FullAdder_364_io_co)
  );
  FullAdder FullAdder_365 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_365_io_a),
    .io_b(FullAdder_365_io_b),
    .io_ci(FullAdder_365_io_ci),
    .io_s(FullAdder_365_io_s),
    .io_co(FullAdder_365_io_co)
  );
  FullAdder FullAdder_366 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_366_io_a),
    .io_b(FullAdder_366_io_b),
    .io_ci(FullAdder_366_io_ci),
    .io_s(FullAdder_366_io_s),
    .io_co(FullAdder_366_io_co)
  );
  FullAdder FullAdder_367 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_367_io_a),
    .io_b(FullAdder_367_io_b),
    .io_ci(FullAdder_367_io_ci),
    .io_s(FullAdder_367_io_s),
    .io_co(FullAdder_367_io_co)
  );
  FullAdder FullAdder_368 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_368_io_a),
    .io_b(FullAdder_368_io_b),
    .io_ci(FullAdder_368_io_ci),
    .io_s(FullAdder_368_io_s),
    .io_co(FullAdder_368_io_co)
  );
  FullAdder FullAdder_369 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_369_io_a),
    .io_b(FullAdder_369_io_b),
    .io_ci(FullAdder_369_io_ci),
    .io_s(FullAdder_369_io_s),
    .io_co(FullAdder_369_io_co)
  );
  FullAdder FullAdder_370 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_370_io_a),
    .io_b(FullAdder_370_io_b),
    .io_ci(FullAdder_370_io_ci),
    .io_s(FullAdder_370_io_s),
    .io_co(FullAdder_370_io_co)
  );
  FullAdder FullAdder_371 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_371_io_a),
    .io_b(FullAdder_371_io_b),
    .io_ci(FullAdder_371_io_ci),
    .io_s(FullAdder_371_io_s),
    .io_co(FullAdder_371_io_co)
  );
  FullAdder FullAdder_372 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_372_io_a),
    .io_b(FullAdder_372_io_b),
    .io_ci(FullAdder_372_io_ci),
    .io_s(FullAdder_372_io_s),
    .io_co(FullAdder_372_io_co)
  );
  FullAdder FullAdder_373 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_373_io_a),
    .io_b(FullAdder_373_io_b),
    .io_ci(FullAdder_373_io_ci),
    .io_s(FullAdder_373_io_s),
    .io_co(FullAdder_373_io_co)
  );
  FullAdder FullAdder_374 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_374_io_a),
    .io_b(FullAdder_374_io_b),
    .io_ci(FullAdder_374_io_ci),
    .io_s(FullAdder_374_io_s),
    .io_co(FullAdder_374_io_co)
  );
  FullAdder FullAdder_375 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_375_io_a),
    .io_b(FullAdder_375_io_b),
    .io_ci(FullAdder_375_io_ci),
    .io_s(FullAdder_375_io_s),
    .io_co(FullAdder_375_io_co)
  );
  FullAdder FullAdder_376 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_376_io_a),
    .io_b(FullAdder_376_io_b),
    .io_ci(FullAdder_376_io_ci),
    .io_s(FullAdder_376_io_s),
    .io_co(FullAdder_376_io_co)
  );
  FullAdder FullAdder_377 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_377_io_a),
    .io_b(FullAdder_377_io_b),
    .io_ci(FullAdder_377_io_ci),
    .io_s(FullAdder_377_io_s),
    .io_co(FullAdder_377_io_co)
  );
  FullAdder FullAdder_378 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_378_io_a),
    .io_b(FullAdder_378_io_b),
    .io_ci(FullAdder_378_io_ci),
    .io_s(FullAdder_378_io_s),
    .io_co(FullAdder_378_io_co)
  );
  HalfAdder HalfAdder_7 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_7_io_a),
    .io_b(HalfAdder_7_io_b),
    .io_s(HalfAdder_7_io_s),
    .io_co(HalfAdder_7_io_co)
  );
  FullAdder FullAdder_379 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_379_io_a),
    .io_b(FullAdder_379_io_b),
    .io_ci(FullAdder_379_io_ci),
    .io_s(FullAdder_379_io_s),
    .io_co(FullAdder_379_io_co)
  );
  FullAdder FullAdder_380 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_380_io_a),
    .io_b(FullAdder_380_io_b),
    .io_ci(FullAdder_380_io_ci),
    .io_s(FullAdder_380_io_s),
    .io_co(FullAdder_380_io_co)
  );
  FullAdder FullAdder_381 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_381_io_a),
    .io_b(FullAdder_381_io_b),
    .io_ci(FullAdder_381_io_ci),
    .io_s(FullAdder_381_io_s),
    .io_co(FullAdder_381_io_co)
  );
  FullAdder FullAdder_382 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_382_io_a),
    .io_b(FullAdder_382_io_b),
    .io_ci(FullAdder_382_io_ci),
    .io_s(FullAdder_382_io_s),
    .io_co(FullAdder_382_io_co)
  );
  FullAdder FullAdder_383 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_383_io_a),
    .io_b(FullAdder_383_io_b),
    .io_ci(FullAdder_383_io_ci),
    .io_s(FullAdder_383_io_s),
    .io_co(FullAdder_383_io_co)
  );
  FullAdder FullAdder_384 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_384_io_a),
    .io_b(FullAdder_384_io_b),
    .io_ci(FullAdder_384_io_ci),
    .io_s(FullAdder_384_io_s),
    .io_co(FullAdder_384_io_co)
  );
  FullAdder FullAdder_385 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_385_io_a),
    .io_b(FullAdder_385_io_b),
    .io_ci(FullAdder_385_io_ci),
    .io_s(FullAdder_385_io_s),
    .io_co(FullAdder_385_io_co)
  );
  FullAdder FullAdder_386 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_386_io_a),
    .io_b(FullAdder_386_io_b),
    .io_ci(FullAdder_386_io_ci),
    .io_s(FullAdder_386_io_s),
    .io_co(FullAdder_386_io_co)
  );
  FullAdder FullAdder_387 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_387_io_a),
    .io_b(FullAdder_387_io_b),
    .io_ci(FullAdder_387_io_ci),
    .io_s(FullAdder_387_io_s),
    .io_co(FullAdder_387_io_co)
  );
  FullAdder FullAdder_388 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_388_io_a),
    .io_b(FullAdder_388_io_b),
    .io_ci(FullAdder_388_io_ci),
    .io_s(FullAdder_388_io_s),
    .io_co(FullAdder_388_io_co)
  );
  FullAdder FullAdder_389 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_389_io_a),
    .io_b(FullAdder_389_io_b),
    .io_ci(FullAdder_389_io_ci),
    .io_s(FullAdder_389_io_s),
    .io_co(FullAdder_389_io_co)
  );
  FullAdder FullAdder_390 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_390_io_a),
    .io_b(FullAdder_390_io_b),
    .io_ci(FullAdder_390_io_ci),
    .io_s(FullAdder_390_io_s),
    .io_co(FullAdder_390_io_co)
  );
  FullAdder FullAdder_391 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_391_io_a),
    .io_b(FullAdder_391_io_b),
    .io_ci(FullAdder_391_io_ci),
    .io_s(FullAdder_391_io_s),
    .io_co(FullAdder_391_io_co)
  );
  HalfAdder HalfAdder_8 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_8_io_a),
    .io_b(HalfAdder_8_io_b),
    .io_s(HalfAdder_8_io_s),
    .io_co(HalfAdder_8_io_co)
  );
  FullAdder FullAdder_392 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_392_io_a),
    .io_b(FullAdder_392_io_b),
    .io_ci(FullAdder_392_io_ci),
    .io_s(FullAdder_392_io_s),
    .io_co(FullAdder_392_io_co)
  );
  FullAdder FullAdder_393 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_393_io_a),
    .io_b(FullAdder_393_io_b),
    .io_ci(FullAdder_393_io_ci),
    .io_s(FullAdder_393_io_s),
    .io_co(FullAdder_393_io_co)
  );
  FullAdder FullAdder_394 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_394_io_a),
    .io_b(FullAdder_394_io_b),
    .io_ci(FullAdder_394_io_ci),
    .io_s(FullAdder_394_io_s),
    .io_co(FullAdder_394_io_co)
  );
  FullAdder FullAdder_395 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_395_io_a),
    .io_b(FullAdder_395_io_b),
    .io_ci(FullAdder_395_io_ci),
    .io_s(FullAdder_395_io_s),
    .io_co(FullAdder_395_io_co)
  );
  FullAdder FullAdder_396 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_396_io_a),
    .io_b(FullAdder_396_io_b),
    .io_ci(FullAdder_396_io_ci),
    .io_s(FullAdder_396_io_s),
    .io_co(FullAdder_396_io_co)
  );
  FullAdder FullAdder_397 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_397_io_a),
    .io_b(FullAdder_397_io_b),
    .io_ci(FullAdder_397_io_ci),
    .io_s(FullAdder_397_io_s),
    .io_co(FullAdder_397_io_co)
  );
  FullAdder FullAdder_398 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_398_io_a),
    .io_b(FullAdder_398_io_b),
    .io_ci(FullAdder_398_io_ci),
    .io_s(FullAdder_398_io_s),
    .io_co(FullAdder_398_io_co)
  );
  FullAdder FullAdder_399 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_399_io_a),
    .io_b(FullAdder_399_io_b),
    .io_ci(FullAdder_399_io_ci),
    .io_s(FullAdder_399_io_s),
    .io_co(FullAdder_399_io_co)
  );
  FullAdder FullAdder_400 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_400_io_a),
    .io_b(FullAdder_400_io_b),
    .io_ci(FullAdder_400_io_ci),
    .io_s(FullAdder_400_io_s),
    .io_co(FullAdder_400_io_co)
  );
  FullAdder FullAdder_401 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_401_io_a),
    .io_b(FullAdder_401_io_b),
    .io_ci(FullAdder_401_io_ci),
    .io_s(FullAdder_401_io_s),
    .io_co(FullAdder_401_io_co)
  );
  FullAdder FullAdder_402 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_402_io_a),
    .io_b(FullAdder_402_io_b),
    .io_ci(FullAdder_402_io_ci),
    .io_s(FullAdder_402_io_s),
    .io_co(FullAdder_402_io_co)
  );
  FullAdder FullAdder_403 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_403_io_a),
    .io_b(FullAdder_403_io_b),
    .io_ci(FullAdder_403_io_ci),
    .io_s(FullAdder_403_io_s),
    .io_co(FullAdder_403_io_co)
  );
  FullAdder FullAdder_404 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_404_io_a),
    .io_b(FullAdder_404_io_b),
    .io_ci(FullAdder_404_io_ci),
    .io_s(FullAdder_404_io_s),
    .io_co(FullAdder_404_io_co)
  );
  HalfAdder HalfAdder_9 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_9_io_a),
    .io_b(HalfAdder_9_io_b),
    .io_s(HalfAdder_9_io_s),
    .io_co(HalfAdder_9_io_co)
  );
  HalfAdder HalfAdder_10 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_10_io_a),
    .io_b(HalfAdder_10_io_b),
    .io_s(HalfAdder_10_io_s),
    .io_co(HalfAdder_10_io_co)
  );
  HalfAdder HalfAdder_11 ( // @[wallaced.scala 77:25]
    .io_a(HalfAdder_11_io_a),
    .io_b(HalfAdder_11_io_b),
    .io_s(HalfAdder_11_io_s),
    .io_co(HalfAdder_11_io_co)
  );
  FullAdder FullAdder_405 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_405_io_a),
    .io_b(FullAdder_405_io_b),
    .io_ci(FullAdder_405_io_ci),
    .io_s(FullAdder_405_io_s),
    .io_co(FullAdder_405_io_co)
  );
  FullAdder FullAdder_406 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_406_io_a),
    .io_b(FullAdder_406_io_b),
    .io_ci(FullAdder_406_io_ci),
    .io_s(FullAdder_406_io_s),
    .io_co(FullAdder_406_io_co)
  );
  FullAdder FullAdder_407 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_407_io_a),
    .io_b(FullAdder_407_io_b),
    .io_ci(FullAdder_407_io_ci),
    .io_s(FullAdder_407_io_s),
    .io_co(FullAdder_407_io_co)
  );
  FullAdder FullAdder_408 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_408_io_a),
    .io_b(FullAdder_408_io_b),
    .io_ci(FullAdder_408_io_ci),
    .io_s(FullAdder_408_io_s),
    .io_co(FullAdder_408_io_co)
  );
  FullAdder FullAdder_409 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_409_io_a),
    .io_b(FullAdder_409_io_b),
    .io_ci(FullAdder_409_io_ci),
    .io_s(FullAdder_409_io_s),
    .io_co(FullAdder_409_io_co)
  );
  FullAdder FullAdder_410 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_410_io_a),
    .io_b(FullAdder_410_io_b),
    .io_ci(FullAdder_410_io_ci),
    .io_s(FullAdder_410_io_s),
    .io_co(FullAdder_410_io_co)
  );
  FullAdder FullAdder_411 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_411_io_a),
    .io_b(FullAdder_411_io_b),
    .io_ci(FullAdder_411_io_ci),
    .io_s(FullAdder_411_io_s),
    .io_co(FullAdder_411_io_co)
  );
  FullAdder FullAdder_412 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_412_io_a),
    .io_b(FullAdder_412_io_b),
    .io_ci(FullAdder_412_io_ci),
    .io_s(FullAdder_412_io_s),
    .io_co(FullAdder_412_io_co)
  );
  FullAdder FullAdder_413 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_413_io_a),
    .io_b(FullAdder_413_io_b),
    .io_ci(FullAdder_413_io_ci),
    .io_s(FullAdder_413_io_s),
    .io_co(FullAdder_413_io_co)
  );
  FullAdder FullAdder_414 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_414_io_a),
    .io_b(FullAdder_414_io_b),
    .io_ci(FullAdder_414_io_ci),
    .io_s(FullAdder_414_io_s),
    .io_co(FullAdder_414_io_co)
  );
  FullAdder FullAdder_415 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_415_io_a),
    .io_b(FullAdder_415_io_b),
    .io_ci(FullAdder_415_io_ci),
    .io_s(FullAdder_415_io_s),
    .io_co(FullAdder_415_io_co)
  );
  FullAdder FullAdder_416 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_416_io_a),
    .io_b(FullAdder_416_io_b),
    .io_ci(FullAdder_416_io_ci),
    .io_s(FullAdder_416_io_s),
    .io_co(FullAdder_416_io_co)
  );
  FullAdder FullAdder_417 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_417_io_a),
    .io_b(FullAdder_417_io_b),
    .io_ci(FullAdder_417_io_ci),
    .io_s(FullAdder_417_io_s),
    .io_co(FullAdder_417_io_co)
  );
  FullAdder FullAdder_418 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_418_io_a),
    .io_b(FullAdder_418_io_b),
    .io_ci(FullAdder_418_io_ci),
    .io_s(FullAdder_418_io_s),
    .io_co(FullAdder_418_io_co)
  );
  FullAdder FullAdder_419 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_419_io_a),
    .io_b(FullAdder_419_io_b),
    .io_ci(FullAdder_419_io_ci),
    .io_s(FullAdder_419_io_s),
    .io_co(FullAdder_419_io_co)
  );
  FullAdder FullAdder_420 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_420_io_a),
    .io_b(FullAdder_420_io_b),
    .io_ci(FullAdder_420_io_ci),
    .io_s(FullAdder_420_io_s),
    .io_co(FullAdder_420_io_co)
  );
  FullAdder FullAdder_421 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_421_io_a),
    .io_b(FullAdder_421_io_b),
    .io_ci(FullAdder_421_io_ci),
    .io_s(FullAdder_421_io_s),
    .io_co(FullAdder_421_io_co)
  );
  FullAdder FullAdder_422 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_422_io_a),
    .io_b(FullAdder_422_io_b),
    .io_ci(FullAdder_422_io_ci),
    .io_s(FullAdder_422_io_s),
    .io_co(FullAdder_422_io_co)
  );
  FullAdder FullAdder_423 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_423_io_a),
    .io_b(FullAdder_423_io_b),
    .io_ci(FullAdder_423_io_ci),
    .io_s(FullAdder_423_io_s),
    .io_co(FullAdder_423_io_co)
  );
  FullAdder FullAdder_424 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_424_io_a),
    .io_b(FullAdder_424_io_b),
    .io_ci(FullAdder_424_io_ci),
    .io_s(FullAdder_424_io_s),
    .io_co(FullAdder_424_io_co)
  );
  FullAdder FullAdder_425 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_425_io_a),
    .io_b(FullAdder_425_io_b),
    .io_ci(FullAdder_425_io_ci),
    .io_s(FullAdder_425_io_s),
    .io_co(FullAdder_425_io_co)
  );
  FullAdder FullAdder_426 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_426_io_a),
    .io_b(FullAdder_426_io_b),
    .io_ci(FullAdder_426_io_ci),
    .io_s(FullAdder_426_io_s),
    .io_co(FullAdder_426_io_co)
  );
  FullAdder FullAdder_427 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_427_io_a),
    .io_b(FullAdder_427_io_b),
    .io_ci(FullAdder_427_io_ci),
    .io_s(FullAdder_427_io_s),
    .io_co(FullAdder_427_io_co)
  );
  FullAdder FullAdder_428 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_428_io_a),
    .io_b(FullAdder_428_io_b),
    .io_ci(FullAdder_428_io_ci),
    .io_s(FullAdder_428_io_s),
    .io_co(FullAdder_428_io_co)
  );
  FullAdder FullAdder_429 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_429_io_a),
    .io_b(FullAdder_429_io_b),
    .io_ci(FullAdder_429_io_ci),
    .io_s(FullAdder_429_io_s),
    .io_co(FullAdder_429_io_co)
  );
  FullAdder FullAdder_430 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_430_io_a),
    .io_b(FullAdder_430_io_b),
    .io_ci(FullAdder_430_io_ci),
    .io_s(FullAdder_430_io_s),
    .io_co(FullAdder_430_io_co)
  );
  FullAdder FullAdder_431 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_431_io_a),
    .io_b(FullAdder_431_io_b),
    .io_ci(FullAdder_431_io_ci),
    .io_s(FullAdder_431_io_s),
    .io_co(FullAdder_431_io_co)
  );
  FullAdder FullAdder_432 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_432_io_a),
    .io_b(FullAdder_432_io_b),
    .io_ci(FullAdder_432_io_ci),
    .io_s(FullAdder_432_io_s),
    .io_co(FullAdder_432_io_co)
  );
  FullAdder FullAdder_433 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_433_io_a),
    .io_b(FullAdder_433_io_b),
    .io_ci(FullAdder_433_io_ci),
    .io_s(FullAdder_433_io_s),
    .io_co(FullAdder_433_io_co)
  );
  FullAdder FullAdder_434 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_434_io_a),
    .io_b(FullAdder_434_io_b),
    .io_ci(FullAdder_434_io_ci),
    .io_s(FullAdder_434_io_s),
    .io_co(FullAdder_434_io_co)
  );
  FullAdder FullAdder_435 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_435_io_a),
    .io_b(FullAdder_435_io_b),
    .io_ci(FullAdder_435_io_ci),
    .io_s(FullAdder_435_io_s),
    .io_co(FullAdder_435_io_co)
  );
  FullAdder FullAdder_436 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_436_io_a),
    .io_b(FullAdder_436_io_b),
    .io_ci(FullAdder_436_io_ci),
    .io_s(FullAdder_436_io_s),
    .io_co(FullAdder_436_io_co)
  );
  FullAdder FullAdder_437 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_437_io_a),
    .io_b(FullAdder_437_io_b),
    .io_ci(FullAdder_437_io_ci),
    .io_s(FullAdder_437_io_s),
    .io_co(FullAdder_437_io_co)
  );
  FullAdder FullAdder_438 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_438_io_a),
    .io_b(FullAdder_438_io_b),
    .io_ci(FullAdder_438_io_ci),
    .io_s(FullAdder_438_io_s),
    .io_co(FullAdder_438_io_co)
  );
  FullAdder FullAdder_439 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_439_io_a),
    .io_b(FullAdder_439_io_b),
    .io_ci(FullAdder_439_io_ci),
    .io_s(FullAdder_439_io_s),
    .io_co(FullAdder_439_io_co)
  );
  FullAdder FullAdder_440 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_440_io_a),
    .io_b(FullAdder_440_io_b),
    .io_ci(FullAdder_440_io_ci),
    .io_s(FullAdder_440_io_s),
    .io_co(FullAdder_440_io_co)
  );
  FullAdder FullAdder_441 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_441_io_a),
    .io_b(FullAdder_441_io_b),
    .io_ci(FullAdder_441_io_ci),
    .io_s(FullAdder_441_io_s),
    .io_co(FullAdder_441_io_co)
  );
  FullAdder FullAdder_442 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_442_io_a),
    .io_b(FullAdder_442_io_b),
    .io_ci(FullAdder_442_io_ci),
    .io_s(FullAdder_442_io_s),
    .io_co(FullAdder_442_io_co)
  );
  FullAdder FullAdder_443 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_443_io_a),
    .io_b(FullAdder_443_io_b),
    .io_ci(FullAdder_443_io_ci),
    .io_s(FullAdder_443_io_s),
    .io_co(FullAdder_443_io_co)
  );
  FullAdder FullAdder_444 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_444_io_a),
    .io_b(FullAdder_444_io_b),
    .io_ci(FullAdder_444_io_ci),
    .io_s(FullAdder_444_io_s),
    .io_co(FullAdder_444_io_co)
  );
  FullAdder FullAdder_445 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_445_io_a),
    .io_b(FullAdder_445_io_b),
    .io_ci(FullAdder_445_io_ci),
    .io_s(FullAdder_445_io_s),
    .io_co(FullAdder_445_io_co)
  );
  FullAdder FullAdder_446 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_446_io_a),
    .io_b(FullAdder_446_io_b),
    .io_ci(FullAdder_446_io_ci),
    .io_s(FullAdder_446_io_s),
    .io_co(FullAdder_446_io_co)
  );
  FullAdder FullAdder_447 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_447_io_a),
    .io_b(FullAdder_447_io_b),
    .io_ci(FullAdder_447_io_ci),
    .io_s(FullAdder_447_io_s),
    .io_co(FullAdder_447_io_co)
  );
  FullAdder FullAdder_448 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_448_io_a),
    .io_b(FullAdder_448_io_b),
    .io_ci(FullAdder_448_io_ci),
    .io_s(FullAdder_448_io_s),
    .io_co(FullAdder_448_io_co)
  );
  FullAdder FullAdder_449 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_449_io_a),
    .io_b(FullAdder_449_io_b),
    .io_ci(FullAdder_449_io_ci),
    .io_s(FullAdder_449_io_s),
    .io_co(FullAdder_449_io_co)
  );
  FullAdder FullAdder_450 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_450_io_a),
    .io_b(FullAdder_450_io_b),
    .io_ci(FullAdder_450_io_ci),
    .io_s(FullAdder_450_io_s),
    .io_co(FullAdder_450_io_co)
  );
  FullAdder FullAdder_451 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_451_io_a),
    .io_b(FullAdder_451_io_b),
    .io_ci(FullAdder_451_io_ci),
    .io_s(FullAdder_451_io_s),
    .io_co(FullAdder_451_io_co)
  );
  FullAdder FullAdder_452 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_452_io_a),
    .io_b(FullAdder_452_io_b),
    .io_ci(FullAdder_452_io_ci),
    .io_s(FullAdder_452_io_s),
    .io_co(FullAdder_452_io_co)
  );
  FullAdder FullAdder_453 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_453_io_a),
    .io_b(FullAdder_453_io_b),
    .io_ci(FullAdder_453_io_ci),
    .io_s(FullAdder_453_io_s),
    .io_co(FullAdder_453_io_co)
  );
  FullAdder FullAdder_454 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_454_io_a),
    .io_b(FullAdder_454_io_b),
    .io_ci(FullAdder_454_io_ci),
    .io_s(FullAdder_454_io_s),
    .io_co(FullAdder_454_io_co)
  );
  FullAdder FullAdder_455 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_455_io_a),
    .io_b(FullAdder_455_io_b),
    .io_ci(FullAdder_455_io_ci),
    .io_s(FullAdder_455_io_s),
    .io_co(FullAdder_455_io_co)
  );
  FullAdder FullAdder_456 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_456_io_a),
    .io_b(FullAdder_456_io_b),
    .io_ci(FullAdder_456_io_ci),
    .io_s(FullAdder_456_io_s),
    .io_co(FullAdder_456_io_co)
  );
  FullAdder FullAdder_457 ( // @[wallaced.scala 86:25]
    .io_a(FullAdder_457_io_a),
    .io_b(FullAdder_457_io_b),
    .io_ci(FullAdder_457_io_ci),
    .io_s(FullAdder_457_io_s),
    .io_co(FullAdder_457_io_co)
  );
  assign io_augend = {_T_541,res0_0}; // @[wallaced.scala 109:13]
  assign io_addend = {_T_572,res1_0}; // @[wallaced.scala 110:13]
  assign FullAdder_io_a = io_pp_13[15]; // @[wallaced.scala 88:18]
  assign FullAdder_io_b = io_pp_14[14]; // @[wallaced.scala 89:18]
  assign FullAdder_io_ci = io_pp_15[13]; // @[wallaced.scala 90:19]
  assign FullAdder_1_io_a = io_pp_12[15]; // @[wallaced.scala 88:18]
  assign FullAdder_1_io_b = io_pp_13[14]; // @[wallaced.scala 89:18]
  assign FullAdder_1_io_ci = io_pp_14[13]; // @[wallaced.scala 90:19]
  assign FullAdder_2_io_a = io_pp_11[15]; // @[wallaced.scala 88:18]
  assign FullAdder_2_io_b = io_pp_12[14]; // @[wallaced.scala 89:18]
  assign FullAdder_2_io_ci = io_pp_13[13]; // @[wallaced.scala 90:19]
  assign FullAdder_3_io_a = io_pp_10[15]; // @[wallaced.scala 88:18]
  assign FullAdder_3_io_b = io_pp_11[14]; // @[wallaced.scala 89:18]
  assign FullAdder_3_io_ci = io_pp_12[13]; // @[wallaced.scala 90:19]
  assign FullAdder_4_io_a = io_pp_13[12]; // @[wallaced.scala 88:18]
  assign FullAdder_4_io_b = io_pp_14[11]; // @[wallaced.scala 89:18]
  assign FullAdder_4_io_ci = io_pp_15[10]; // @[wallaced.scala 90:19]
  assign FullAdder_5_io_a = io_pp_9[15]; // @[wallaced.scala 88:18]
  assign FullAdder_5_io_b = io_pp_10[14]; // @[wallaced.scala 89:18]
  assign FullAdder_5_io_ci = io_pp_11[13]; // @[wallaced.scala 90:19]
  assign FullAdder_6_io_a = io_pp_12[12]; // @[wallaced.scala 88:18]
  assign FullAdder_6_io_b = io_pp_13[11]; // @[wallaced.scala 89:18]
  assign FullAdder_6_io_ci = io_pp_14[10]; // @[wallaced.scala 90:19]
  assign FullAdder_7_io_a = io_pp_8[15]; // @[wallaced.scala 88:18]
  assign FullAdder_7_io_b = io_pp_9[14]; // @[wallaced.scala 89:18]
  assign FullAdder_7_io_ci = io_pp_10[13]; // @[wallaced.scala 90:19]
  assign FullAdder_8_io_a = io_pp_11[12]; // @[wallaced.scala 88:18]
  assign FullAdder_8_io_b = io_pp_12[11]; // @[wallaced.scala 89:18]
  assign FullAdder_8_io_ci = io_pp_13[10]; // @[wallaced.scala 90:19]
  assign FullAdder_9_io_a = io_pp_7[15]; // @[wallaced.scala 88:18]
  assign FullAdder_9_io_b = io_pp_8[14]; // @[wallaced.scala 89:18]
  assign FullAdder_9_io_ci = io_pp_9[13]; // @[wallaced.scala 90:19]
  assign FullAdder_10_io_a = io_pp_10[12]; // @[wallaced.scala 88:18]
  assign FullAdder_10_io_b = io_pp_11[11]; // @[wallaced.scala 89:18]
  assign FullAdder_10_io_ci = io_pp_12[10]; // @[wallaced.scala 90:19]
  assign FullAdder_11_io_a = io_pp_13[9]; // @[wallaced.scala 88:18]
  assign FullAdder_11_io_b = io_pp_14[8]; // @[wallaced.scala 89:18]
  assign FullAdder_11_io_ci = io_pp_15[7]; // @[wallaced.scala 90:19]
  assign FullAdder_12_io_a = io_pp_6[15]; // @[wallaced.scala 88:18]
  assign FullAdder_12_io_b = io_pp_7[14]; // @[wallaced.scala 89:18]
  assign FullAdder_12_io_ci = io_pp_8[13]; // @[wallaced.scala 90:19]
  assign FullAdder_13_io_a = io_pp_9[12]; // @[wallaced.scala 88:18]
  assign FullAdder_13_io_b = io_pp_10[11]; // @[wallaced.scala 89:18]
  assign FullAdder_13_io_ci = io_pp_11[10]; // @[wallaced.scala 90:19]
  assign FullAdder_14_io_a = io_pp_12[9]; // @[wallaced.scala 88:18]
  assign FullAdder_14_io_b = io_pp_13[8]; // @[wallaced.scala 89:18]
  assign FullAdder_14_io_ci = io_pp_14[7]; // @[wallaced.scala 90:19]
  assign FullAdder_15_io_a = io_pp_5[15]; // @[wallaced.scala 88:18]
  assign FullAdder_15_io_b = io_pp_6[14]; // @[wallaced.scala 89:18]
  assign FullAdder_15_io_ci = io_pp_7[13]; // @[wallaced.scala 90:19]
  assign FullAdder_16_io_a = io_pp_8[12]; // @[wallaced.scala 88:18]
  assign FullAdder_16_io_b = io_pp_9[11]; // @[wallaced.scala 89:18]
  assign FullAdder_16_io_ci = io_pp_10[10]; // @[wallaced.scala 90:19]
  assign FullAdder_17_io_a = io_pp_11[9]; // @[wallaced.scala 88:18]
  assign FullAdder_17_io_b = io_pp_12[8]; // @[wallaced.scala 89:18]
  assign FullAdder_17_io_ci = io_pp_13[7]; // @[wallaced.scala 90:19]
  assign FullAdder_18_io_a = io_pp_4[15]; // @[wallaced.scala 88:18]
  assign FullAdder_18_io_b = io_pp_5[14]; // @[wallaced.scala 89:18]
  assign FullAdder_18_io_ci = io_pp_6[13]; // @[wallaced.scala 90:19]
  assign FullAdder_19_io_a = io_pp_7[12]; // @[wallaced.scala 88:18]
  assign FullAdder_19_io_b = io_pp_8[11]; // @[wallaced.scala 89:18]
  assign FullAdder_19_io_ci = io_pp_9[10]; // @[wallaced.scala 90:19]
  assign FullAdder_20_io_a = io_pp_10[9]; // @[wallaced.scala 88:18]
  assign FullAdder_20_io_b = io_pp_11[8]; // @[wallaced.scala 89:18]
  assign FullAdder_20_io_ci = io_pp_12[7]; // @[wallaced.scala 90:19]
  assign FullAdder_21_io_a = io_pp_13[6]; // @[wallaced.scala 88:18]
  assign FullAdder_21_io_b = io_pp_14[5]; // @[wallaced.scala 89:18]
  assign FullAdder_21_io_ci = io_pp_15[4]; // @[wallaced.scala 90:19]
  assign FullAdder_22_io_a = io_pp_3[15]; // @[wallaced.scala 88:18]
  assign FullAdder_22_io_b = io_pp_4[14]; // @[wallaced.scala 89:18]
  assign FullAdder_22_io_ci = io_pp_5[13]; // @[wallaced.scala 90:19]
  assign FullAdder_23_io_a = io_pp_6[12]; // @[wallaced.scala 88:18]
  assign FullAdder_23_io_b = io_pp_7[11]; // @[wallaced.scala 89:18]
  assign FullAdder_23_io_ci = io_pp_8[10]; // @[wallaced.scala 90:19]
  assign FullAdder_24_io_a = io_pp_9[9]; // @[wallaced.scala 88:18]
  assign FullAdder_24_io_b = io_pp_10[8]; // @[wallaced.scala 89:18]
  assign FullAdder_24_io_ci = io_pp_11[7]; // @[wallaced.scala 90:19]
  assign FullAdder_25_io_a = io_pp_12[6]; // @[wallaced.scala 88:18]
  assign FullAdder_25_io_b = io_pp_13[5]; // @[wallaced.scala 89:18]
  assign FullAdder_25_io_ci = io_pp_14[4]; // @[wallaced.scala 90:19]
  assign FullAdder_26_io_a = io_pp_2[15]; // @[wallaced.scala 88:18]
  assign FullAdder_26_io_b = io_pp_3[14]; // @[wallaced.scala 89:18]
  assign FullAdder_26_io_ci = io_pp_4[13]; // @[wallaced.scala 90:19]
  assign FullAdder_27_io_a = io_pp_5[12]; // @[wallaced.scala 88:18]
  assign FullAdder_27_io_b = io_pp_6[11]; // @[wallaced.scala 89:18]
  assign FullAdder_27_io_ci = io_pp_7[10]; // @[wallaced.scala 90:19]
  assign FullAdder_28_io_a = io_pp_8[9]; // @[wallaced.scala 88:18]
  assign FullAdder_28_io_b = io_pp_9[8]; // @[wallaced.scala 89:18]
  assign FullAdder_28_io_ci = io_pp_10[7]; // @[wallaced.scala 90:19]
  assign FullAdder_29_io_a = io_pp_11[6]; // @[wallaced.scala 88:18]
  assign FullAdder_29_io_b = io_pp_12[5]; // @[wallaced.scala 89:18]
  assign FullAdder_29_io_ci = io_pp_13[4]; // @[wallaced.scala 90:19]
  assign FullAdder_30_io_a = io_pp_1[15]; // @[wallaced.scala 88:18]
  assign FullAdder_30_io_b = io_pp_2[14]; // @[wallaced.scala 89:18]
  assign FullAdder_30_io_ci = io_pp_3[13]; // @[wallaced.scala 90:19]
  assign FullAdder_31_io_a = io_pp_4[12]; // @[wallaced.scala 88:18]
  assign FullAdder_31_io_b = io_pp_5[11]; // @[wallaced.scala 89:18]
  assign FullAdder_31_io_ci = io_pp_6[10]; // @[wallaced.scala 90:19]
  assign FullAdder_32_io_a = io_pp_7[9]; // @[wallaced.scala 88:18]
  assign FullAdder_32_io_b = io_pp_8[8]; // @[wallaced.scala 89:18]
  assign FullAdder_32_io_ci = io_pp_9[7]; // @[wallaced.scala 90:19]
  assign FullAdder_33_io_a = io_pp_10[6]; // @[wallaced.scala 88:18]
  assign FullAdder_33_io_b = io_pp_11[5]; // @[wallaced.scala 89:18]
  assign FullAdder_33_io_ci = io_pp_12[4]; // @[wallaced.scala 90:19]
  assign FullAdder_34_io_a = io_pp_13[3]; // @[wallaced.scala 88:18]
  assign FullAdder_34_io_b = io_pp_14[2]; // @[wallaced.scala 89:18]
  assign FullAdder_34_io_ci = io_pp_15[1]; // @[wallaced.scala 90:19]
  assign FullAdder_35_io_a = io_pp_0[15]; // @[wallaced.scala 88:18]
  assign FullAdder_35_io_b = io_pp_1[14]; // @[wallaced.scala 89:18]
  assign FullAdder_35_io_ci = io_pp_2[13]; // @[wallaced.scala 90:19]
  assign FullAdder_36_io_a = io_pp_3[12]; // @[wallaced.scala 88:18]
  assign FullAdder_36_io_b = io_pp_4[11]; // @[wallaced.scala 89:18]
  assign FullAdder_36_io_ci = io_pp_5[10]; // @[wallaced.scala 90:19]
  assign FullAdder_37_io_a = io_pp_6[9]; // @[wallaced.scala 88:18]
  assign FullAdder_37_io_b = io_pp_7[8]; // @[wallaced.scala 89:18]
  assign FullAdder_37_io_ci = io_pp_8[7]; // @[wallaced.scala 90:19]
  assign FullAdder_38_io_a = io_pp_9[6]; // @[wallaced.scala 88:18]
  assign FullAdder_38_io_b = io_pp_10[5]; // @[wallaced.scala 89:18]
  assign FullAdder_38_io_ci = io_pp_11[4]; // @[wallaced.scala 90:19]
  assign FullAdder_39_io_a = io_pp_12[3]; // @[wallaced.scala 88:18]
  assign FullAdder_39_io_b = io_pp_13[2]; // @[wallaced.scala 89:18]
  assign FullAdder_39_io_ci = io_pp_14[1]; // @[wallaced.scala 90:19]
  assign FullAdder_40_io_a = io_pp_0[14]; // @[wallaced.scala 88:18]
  assign FullAdder_40_io_b = io_pp_1[13]; // @[wallaced.scala 89:18]
  assign FullAdder_40_io_ci = io_pp_2[12]; // @[wallaced.scala 90:19]
  assign FullAdder_41_io_a = io_pp_3[11]; // @[wallaced.scala 88:18]
  assign FullAdder_41_io_b = io_pp_4[10]; // @[wallaced.scala 89:18]
  assign FullAdder_41_io_ci = io_pp_5[9]; // @[wallaced.scala 90:19]
  assign FullAdder_42_io_a = io_pp_6[8]; // @[wallaced.scala 88:18]
  assign FullAdder_42_io_b = io_pp_7[7]; // @[wallaced.scala 89:18]
  assign FullAdder_42_io_ci = io_pp_8[6]; // @[wallaced.scala 90:19]
  assign FullAdder_43_io_a = io_pp_9[5]; // @[wallaced.scala 88:18]
  assign FullAdder_43_io_b = io_pp_10[4]; // @[wallaced.scala 89:18]
  assign FullAdder_43_io_ci = io_pp_11[3]; // @[wallaced.scala 90:19]
  assign FullAdder_44_io_a = io_pp_12[2]; // @[wallaced.scala 88:18]
  assign FullAdder_44_io_b = io_pp_13[1]; // @[wallaced.scala 89:18]
  assign FullAdder_44_io_ci = io_pp_14[0]; // @[wallaced.scala 90:19]
  assign FullAdder_45_io_a = io_pp_0[13]; // @[wallaced.scala 88:18]
  assign FullAdder_45_io_b = io_pp_1[12]; // @[wallaced.scala 89:18]
  assign FullAdder_45_io_ci = io_pp_2[11]; // @[wallaced.scala 90:19]
  assign FullAdder_46_io_a = io_pp_3[10]; // @[wallaced.scala 88:18]
  assign FullAdder_46_io_b = io_pp_4[9]; // @[wallaced.scala 89:18]
  assign FullAdder_46_io_ci = io_pp_5[8]; // @[wallaced.scala 90:19]
  assign FullAdder_47_io_a = io_pp_6[7]; // @[wallaced.scala 88:18]
  assign FullAdder_47_io_b = io_pp_7[6]; // @[wallaced.scala 89:18]
  assign FullAdder_47_io_ci = io_pp_8[5]; // @[wallaced.scala 90:19]
  assign FullAdder_48_io_a = io_pp_9[4]; // @[wallaced.scala 88:18]
  assign FullAdder_48_io_b = io_pp_10[3]; // @[wallaced.scala 89:18]
  assign FullAdder_48_io_ci = io_pp_11[2]; // @[wallaced.scala 90:19]
  assign FullAdder_49_io_a = io_pp_0[12]; // @[wallaced.scala 88:18]
  assign FullAdder_49_io_b = io_pp_1[11]; // @[wallaced.scala 89:18]
  assign FullAdder_49_io_ci = io_pp_2[10]; // @[wallaced.scala 90:19]
  assign FullAdder_50_io_a = io_pp_3[9]; // @[wallaced.scala 88:18]
  assign FullAdder_50_io_b = io_pp_4[8]; // @[wallaced.scala 89:18]
  assign FullAdder_50_io_ci = io_pp_5[7]; // @[wallaced.scala 90:19]
  assign FullAdder_51_io_a = io_pp_6[6]; // @[wallaced.scala 88:18]
  assign FullAdder_51_io_b = io_pp_7[5]; // @[wallaced.scala 89:18]
  assign FullAdder_51_io_ci = io_pp_8[4]; // @[wallaced.scala 90:19]
  assign FullAdder_52_io_a = io_pp_9[3]; // @[wallaced.scala 88:18]
  assign FullAdder_52_io_b = io_pp_10[2]; // @[wallaced.scala 89:18]
  assign FullAdder_52_io_ci = io_pp_11[1]; // @[wallaced.scala 90:19]
  assign FullAdder_53_io_a = io_pp_0[11]; // @[wallaced.scala 88:18]
  assign FullAdder_53_io_b = io_pp_1[10]; // @[wallaced.scala 89:18]
  assign FullAdder_53_io_ci = io_pp_2[9]; // @[wallaced.scala 90:19]
  assign FullAdder_54_io_a = io_pp_3[8]; // @[wallaced.scala 88:18]
  assign FullAdder_54_io_b = io_pp_4[7]; // @[wallaced.scala 89:18]
  assign FullAdder_54_io_ci = io_pp_5[6]; // @[wallaced.scala 90:19]
  assign FullAdder_55_io_a = io_pp_6[5]; // @[wallaced.scala 88:18]
  assign FullAdder_55_io_b = io_pp_7[4]; // @[wallaced.scala 89:18]
  assign FullAdder_55_io_ci = io_pp_8[3]; // @[wallaced.scala 90:19]
  assign FullAdder_56_io_a = io_pp_9[2]; // @[wallaced.scala 88:18]
  assign FullAdder_56_io_b = io_pp_10[1]; // @[wallaced.scala 89:18]
  assign FullAdder_56_io_ci = io_pp_11[0]; // @[wallaced.scala 90:19]
  assign FullAdder_57_io_a = io_pp_0[10]; // @[wallaced.scala 88:18]
  assign FullAdder_57_io_b = io_pp_1[9]; // @[wallaced.scala 89:18]
  assign FullAdder_57_io_ci = io_pp_2[8]; // @[wallaced.scala 90:19]
  assign FullAdder_58_io_a = io_pp_3[7]; // @[wallaced.scala 88:18]
  assign FullAdder_58_io_b = io_pp_4[6]; // @[wallaced.scala 89:18]
  assign FullAdder_58_io_ci = io_pp_5[5]; // @[wallaced.scala 90:19]
  assign FullAdder_59_io_a = io_pp_6[4]; // @[wallaced.scala 88:18]
  assign FullAdder_59_io_b = io_pp_7[3]; // @[wallaced.scala 89:18]
  assign FullAdder_59_io_ci = io_pp_8[2]; // @[wallaced.scala 90:19]
  assign FullAdder_60_io_a = io_pp_0[9]; // @[wallaced.scala 88:18]
  assign FullAdder_60_io_b = io_pp_1[8]; // @[wallaced.scala 89:18]
  assign FullAdder_60_io_ci = io_pp_2[7]; // @[wallaced.scala 90:19]
  assign FullAdder_61_io_a = io_pp_3[6]; // @[wallaced.scala 88:18]
  assign FullAdder_61_io_b = io_pp_4[5]; // @[wallaced.scala 89:18]
  assign FullAdder_61_io_ci = io_pp_5[4]; // @[wallaced.scala 90:19]
  assign FullAdder_62_io_a = io_pp_6[3]; // @[wallaced.scala 88:18]
  assign FullAdder_62_io_b = io_pp_7[2]; // @[wallaced.scala 89:18]
  assign FullAdder_62_io_ci = io_pp_8[1]; // @[wallaced.scala 90:19]
  assign FullAdder_63_io_a = io_pp_0[8]; // @[wallaced.scala 88:18]
  assign FullAdder_63_io_b = io_pp_1[7]; // @[wallaced.scala 89:18]
  assign FullAdder_63_io_ci = io_pp_2[6]; // @[wallaced.scala 90:19]
  assign FullAdder_64_io_a = io_pp_3[5]; // @[wallaced.scala 88:18]
  assign FullAdder_64_io_b = io_pp_4[4]; // @[wallaced.scala 89:18]
  assign FullAdder_64_io_ci = io_pp_5[3]; // @[wallaced.scala 90:19]
  assign FullAdder_65_io_a = io_pp_6[2]; // @[wallaced.scala 88:18]
  assign FullAdder_65_io_b = io_pp_7[1]; // @[wallaced.scala 89:18]
  assign FullAdder_65_io_ci = io_pp_8[0]; // @[wallaced.scala 90:19]
  assign FullAdder_66_io_a = io_pp_0[7]; // @[wallaced.scala 88:18]
  assign FullAdder_66_io_b = io_pp_1[6]; // @[wallaced.scala 89:18]
  assign FullAdder_66_io_ci = io_pp_2[5]; // @[wallaced.scala 90:19]
  assign FullAdder_67_io_a = io_pp_3[4]; // @[wallaced.scala 88:18]
  assign FullAdder_67_io_b = io_pp_4[3]; // @[wallaced.scala 89:18]
  assign FullAdder_67_io_ci = io_pp_5[2]; // @[wallaced.scala 90:19]
  assign FullAdder_68_io_a = io_pp_0[6]; // @[wallaced.scala 88:18]
  assign FullAdder_68_io_b = io_pp_1[5]; // @[wallaced.scala 89:18]
  assign FullAdder_68_io_ci = io_pp_2[4]; // @[wallaced.scala 90:19]
  assign FullAdder_69_io_a = io_pp_3[3]; // @[wallaced.scala 88:18]
  assign FullAdder_69_io_b = io_pp_4[2]; // @[wallaced.scala 89:18]
  assign FullAdder_69_io_ci = io_pp_5[1]; // @[wallaced.scala 90:19]
  assign FullAdder_70_io_a = io_pp_0[5]; // @[wallaced.scala 88:18]
  assign FullAdder_70_io_b = io_pp_1[4]; // @[wallaced.scala 89:18]
  assign FullAdder_70_io_ci = io_pp_2[3]; // @[wallaced.scala 90:19]
  assign FullAdder_71_io_a = io_pp_3[2]; // @[wallaced.scala 88:18]
  assign FullAdder_71_io_b = io_pp_4[1]; // @[wallaced.scala 89:18]
  assign FullAdder_71_io_ci = io_pp_5[0]; // @[wallaced.scala 90:19]
  assign FullAdder_72_io_a = io_pp_0[4]; // @[wallaced.scala 88:18]
  assign FullAdder_72_io_b = io_pp_1[3]; // @[wallaced.scala 89:18]
  assign FullAdder_72_io_ci = io_pp_2[2]; // @[wallaced.scala 90:19]
  assign FullAdder_73_io_a = io_pp_0[3]; // @[wallaced.scala 88:18]
  assign FullAdder_73_io_b = io_pp_1[2]; // @[wallaced.scala 89:18]
  assign FullAdder_73_io_ci = io_pp_2[1]; // @[wallaced.scala 90:19]
  assign FullAdder_74_io_a = io_pp_0[2]; // @[wallaced.scala 88:18]
  assign FullAdder_74_io_b = io_pp_1[1]; // @[wallaced.scala 89:18]
  assign FullAdder_74_io_ci = io_pp_2[0]; // @[wallaced.scala 90:19]
  assign FullAdder_75_io_a = io_pp_14[15]; // @[wallaced.scala 88:18]
  assign FullAdder_75_io_b = io_pp_15[14]; // @[wallaced.scala 89:18]
  assign FullAdder_75_io_ci = io_pp_30[15]; // @[wallaced.scala 90:19]
  assign FullAdder_76_io_a = io_pp_15[12]; // @[wallaced.scala 88:18]
  assign FullAdder_76_io_b = io_pp_28[15]; // @[wallaced.scala 89:18]
  assign FullAdder_76_io_ci = io_pp_29[14]; // @[wallaced.scala 90:19]
  assign FullAdder_77_io_a = io_pp_14[12]; // @[wallaced.scala 88:18]
  assign FullAdder_77_io_b = io_pp_15[11]; // @[wallaced.scala 89:18]
  assign FullAdder_77_io_ci = io_pp_27[15]; // @[wallaced.scala 90:19]
  assign FullAdder_78_io_a = io_pp_26[15]; // @[wallaced.scala 88:18]
  assign FullAdder_78_io_b = io_pp_27[14]; // @[wallaced.scala 89:18]
  assign FullAdder_78_io_ci = io_pp_28[13]; // @[wallaced.scala 90:19]
  assign FullAdder_79_io_a = io_pp_15[9]; // @[wallaced.scala 88:18]
  assign FullAdder_79_io_b = io_pp_25[15]; // @[wallaced.scala 89:18]
  assign FullAdder_79_io_ci = io_pp_26[14]; // @[wallaced.scala 90:19]
  assign FullAdder_80_io_a = io_pp_14[9]; // @[wallaced.scala 88:18]
  assign FullAdder_80_io_b = io_pp_15[8]; // @[wallaced.scala 89:18]
  assign FullAdder_80_io_ci = io_pp_24[15]; // @[wallaced.scala 90:19]
  assign FullAdder_81_io_a = io_pp_25[14]; // @[wallaced.scala 88:18]
  assign FullAdder_81_io_b = io_pp_26[13]; // @[wallaced.scala 89:18]
  assign FullAdder_81_io_ci = io_pp_27[12]; // @[wallaced.scala 90:19]
  assign FullAdder_82_io_a = io_pp_23[15]; // @[wallaced.scala 88:18]
  assign FullAdder_82_io_b = io_pp_24[14]; // @[wallaced.scala 89:18]
  assign FullAdder_82_io_ci = io_pp_25[13]; // @[wallaced.scala 90:19]
  assign FullAdder_83_io_a = io_pp_26[12]; // @[wallaced.scala 88:18]
  assign FullAdder_83_io_b = io_pp_27[11]; // @[wallaced.scala 89:18]
  assign FullAdder_83_io_ci = io_pp_28[10]; // @[wallaced.scala 90:19]
  assign FullAdder_84_io_a = io_pp_15[6]; // @[wallaced.scala 88:18]
  assign FullAdder_84_io_b = io_pp_22[15]; // @[wallaced.scala 89:18]
  assign FullAdder_84_io_ci = io_pp_23[14]; // @[wallaced.scala 90:19]
  assign FullAdder_85_io_a = io_pp_24[13]; // @[wallaced.scala 88:18]
  assign FullAdder_85_io_b = io_pp_25[12]; // @[wallaced.scala 89:18]
  assign FullAdder_85_io_ci = io_pp_26[11]; // @[wallaced.scala 90:19]
  assign FullAdder_86_io_a = io_pp_14[6]; // @[wallaced.scala 88:18]
  assign FullAdder_86_io_b = io_pp_15[5]; // @[wallaced.scala 89:18]
  assign FullAdder_86_io_ci = io_pp_21[15]; // @[wallaced.scala 90:19]
  assign FullAdder_87_io_a = io_pp_22[14]; // @[wallaced.scala 88:18]
  assign FullAdder_87_io_b = io_pp_23[13]; // @[wallaced.scala 89:18]
  assign FullAdder_87_io_ci = io_pp_24[12]; // @[wallaced.scala 90:19]
  assign FullAdder_88_io_a = io_pp_25[11]; // @[wallaced.scala 88:18]
  assign FullAdder_88_io_b = io_pp_26[10]; // @[wallaced.scala 89:18]
  assign FullAdder_88_io_ci = io_pp_27[9]; // @[wallaced.scala 90:19]
  assign FullAdder_89_io_a = io_pp_20[15]; // @[wallaced.scala 88:18]
  assign FullAdder_89_io_b = io_pp_21[14]; // @[wallaced.scala 89:18]
  assign FullAdder_89_io_ci = io_pp_22[13]; // @[wallaced.scala 90:19]
  assign FullAdder_90_io_a = io_pp_23[12]; // @[wallaced.scala 88:18]
  assign FullAdder_90_io_b = io_pp_24[11]; // @[wallaced.scala 89:18]
  assign FullAdder_90_io_ci = io_pp_25[10]; // @[wallaced.scala 90:19]
  assign FullAdder_91_io_a = io_pp_15[3]; // @[wallaced.scala 88:18]
  assign FullAdder_91_io_b = io_pp_19[15]; // @[wallaced.scala 89:18]
  assign FullAdder_91_io_ci = io_pp_20[14]; // @[wallaced.scala 90:19]
  assign FullAdder_92_io_a = io_pp_21[13]; // @[wallaced.scala 88:18]
  assign FullAdder_92_io_b = io_pp_22[12]; // @[wallaced.scala 89:18]
  assign FullAdder_92_io_ci = io_pp_23[11]; // @[wallaced.scala 90:19]
  assign FullAdder_93_io_a = io_pp_24[10]; // @[wallaced.scala 88:18]
  assign FullAdder_93_io_b = io_pp_25[9]; // @[wallaced.scala 89:18]
  assign FullAdder_93_io_ci = io_pp_26[8]; // @[wallaced.scala 90:19]
  assign FullAdder_94_io_a = io_pp_14[3]; // @[wallaced.scala 88:18]
  assign FullAdder_94_io_b = io_pp_15[2]; // @[wallaced.scala 89:18]
  assign FullAdder_94_io_ci = io_pp_18[15]; // @[wallaced.scala 90:19]
  assign FullAdder_95_io_a = io_pp_19[14]; // @[wallaced.scala 88:18]
  assign FullAdder_95_io_b = io_pp_20[13]; // @[wallaced.scala 89:18]
  assign FullAdder_95_io_ci = io_pp_21[12]; // @[wallaced.scala 90:19]
  assign FullAdder_96_io_a = io_pp_22[11]; // @[wallaced.scala 88:18]
  assign FullAdder_96_io_b = io_pp_23[10]; // @[wallaced.scala 89:18]
  assign FullAdder_96_io_ci = io_pp_24[9]; // @[wallaced.scala 90:19]
  assign FullAdder_97_io_a = io_pp_17[15]; // @[wallaced.scala 88:18]
  assign FullAdder_97_io_b = io_pp_18[14]; // @[wallaced.scala 89:18]
  assign FullAdder_97_io_ci = io_pp_19[13]; // @[wallaced.scala 90:19]
  assign FullAdder_98_io_a = io_pp_20[12]; // @[wallaced.scala 88:18]
  assign FullAdder_98_io_b = io_pp_21[11]; // @[wallaced.scala 89:18]
  assign FullAdder_98_io_ci = io_pp_22[10]; // @[wallaced.scala 90:19]
  assign FullAdder_99_io_a = io_pp_23[9]; // @[wallaced.scala 88:18]
  assign FullAdder_99_io_b = io_pp_24[8]; // @[wallaced.scala 89:18]
  assign FullAdder_99_io_ci = io_pp_25[7]; // @[wallaced.scala 90:19]
  assign FullAdder_100_io_a = io_pp_15[0]; // @[wallaced.scala 88:18]
  assign FullAdder_100_io_b = io_pp_16[15]; // @[wallaced.scala 89:18]
  assign FullAdder_100_io_ci = io_pp_17[14]; // @[wallaced.scala 90:19]
  assign FullAdder_101_io_a = io_pp_18[13]; // @[wallaced.scala 88:18]
  assign FullAdder_101_io_b = io_pp_19[12]; // @[wallaced.scala 89:18]
  assign FullAdder_101_io_ci = io_pp_20[11]; // @[wallaced.scala 90:19]
  assign FullAdder_102_io_a = io_pp_21[10]; // @[wallaced.scala 88:18]
  assign FullAdder_102_io_b = io_pp_22[9]; // @[wallaced.scala 89:18]
  assign FullAdder_102_io_ci = io_pp_23[8]; // @[wallaced.scala 90:19]
  assign FullAdder_103_io_a = io_pp_16[14]; // @[wallaced.scala 88:18]
  assign FullAdder_103_io_b = io_pp_17[13]; // @[wallaced.scala 89:18]
  assign FullAdder_103_io_ci = io_pp_18[12]; // @[wallaced.scala 90:19]
  assign FullAdder_104_io_a = io_pp_19[11]; // @[wallaced.scala 88:18]
  assign FullAdder_104_io_b = io_pp_20[10]; // @[wallaced.scala 89:18]
  assign FullAdder_104_io_ci = io_pp_21[9]; // @[wallaced.scala 90:19]
  assign FullAdder_105_io_a = io_pp_22[8]; // @[wallaced.scala 88:18]
  assign FullAdder_105_io_b = io_pp_23[7]; // @[wallaced.scala 89:18]
  assign FullAdder_105_io_ci = io_pp_24[6]; // @[wallaced.scala 90:19]
  assign FullAdder_106_io_a = io_pp_12[1]; // @[wallaced.scala 88:18]
  assign FullAdder_106_io_b = io_pp_13[0]; // @[wallaced.scala 89:18]
  assign FullAdder_106_io_ci = io_pp_16[13]; // @[wallaced.scala 90:19]
  assign FullAdder_107_io_a = io_pp_17[12]; // @[wallaced.scala 88:18]
  assign FullAdder_107_io_b = io_pp_18[11]; // @[wallaced.scala 89:18]
  assign FullAdder_107_io_ci = io_pp_19[10]; // @[wallaced.scala 90:19]
  assign FullAdder_108_io_a = io_pp_20[9]; // @[wallaced.scala 88:18]
  assign FullAdder_108_io_b = io_pp_21[8]; // @[wallaced.scala 89:18]
  assign FullAdder_108_io_ci = io_pp_22[7]; // @[wallaced.scala 90:19]
  assign FullAdder_109_io_a = io_pp_12[0]; // @[wallaced.scala 88:18]
  assign FullAdder_109_io_b = io_pp_16[12]; // @[wallaced.scala 89:18]
  assign FullAdder_109_io_ci = io_pp_17[11]; // @[wallaced.scala 90:19]
  assign FullAdder_110_io_a = io_pp_18[10]; // @[wallaced.scala 88:18]
  assign FullAdder_110_io_b = io_pp_19[9]; // @[wallaced.scala 89:18]
  assign FullAdder_110_io_ci = io_pp_20[8]; // @[wallaced.scala 90:19]
  assign FullAdder_111_io_a = io_pp_21[7]; // @[wallaced.scala 88:18]
  assign FullAdder_111_io_b = io_pp_22[6]; // @[wallaced.scala 89:18]
  assign FullAdder_111_io_ci = io_pp_23[5]; // @[wallaced.scala 90:19]
  assign FullAdder_112_io_a = io_pp_16[11]; // @[wallaced.scala 88:18]
  assign FullAdder_112_io_b = io_pp_17[10]; // @[wallaced.scala 89:18]
  assign FullAdder_112_io_ci = io_pp_18[9]; // @[wallaced.scala 90:19]
  assign FullAdder_113_io_a = io_pp_19[8]; // @[wallaced.scala 88:18]
  assign FullAdder_113_io_b = io_pp_20[7]; // @[wallaced.scala 89:18]
  assign FullAdder_113_io_ci = io_pp_21[6]; // @[wallaced.scala 90:19]
  assign FullAdder_114_io_a = io_pp_9[1]; // @[wallaced.scala 88:18]
  assign FullAdder_114_io_b = io_pp_10[0]; // @[wallaced.scala 89:18]
  assign FullAdder_114_io_ci = io_pp_16[10]; // @[wallaced.scala 90:19]
  assign FullAdder_115_io_a = io_pp_17[9]; // @[wallaced.scala 88:18]
  assign FullAdder_115_io_b = io_pp_18[8]; // @[wallaced.scala 89:18]
  assign FullAdder_115_io_ci = io_pp_19[7]; // @[wallaced.scala 90:19]
  assign FullAdder_116_io_a = io_pp_9[0]; // @[wallaced.scala 88:18]
  assign FullAdder_116_io_b = io_pp_16[9]; // @[wallaced.scala 89:18]
  assign FullAdder_116_io_ci = io_pp_17[8]; // @[wallaced.scala 90:19]
  assign FullAdder_117_io_a = io_pp_18[7]; // @[wallaced.scala 88:18]
  assign FullAdder_117_io_b = io_pp_19[6]; // @[wallaced.scala 89:18]
  assign FullAdder_117_io_ci = io_pp_20[5]; // @[wallaced.scala 90:19]
  assign FullAdder_118_io_a = io_pp_16[8]; // @[wallaced.scala 88:18]
  assign FullAdder_118_io_b = io_pp_17[7]; // @[wallaced.scala 89:18]
  assign FullAdder_118_io_ci = io_pp_18[6]; // @[wallaced.scala 90:19]
  assign FullAdder_119_io_a = io_pp_6[1]; // @[wallaced.scala 88:18]
  assign FullAdder_119_io_b = io_pp_7[0]; // @[wallaced.scala 89:18]
  assign FullAdder_119_io_ci = io_pp_16[7]; // @[wallaced.scala 90:19]
  assign FullAdder_120_io_a = io_pp_17[6]; // @[wallaced.scala 88:18]
  assign FullAdder_120_io_b = io_pp_18[5]; // @[wallaced.scala 89:18]
  assign FullAdder_120_io_ci = io_pp_19[4]; // @[wallaced.scala 90:19]
  assign FullAdder_121_io_a = io_pp_6[0]; // @[wallaced.scala 88:18]
  assign FullAdder_121_io_b = io_pp_16[6]; // @[wallaced.scala 89:18]
  assign FullAdder_121_io_ci = io_pp_17[5]; // @[wallaced.scala 90:19]
  assign FullAdder_122_io_a = io_pp_16[5]; // @[wallaced.scala 88:18]
  assign FullAdder_122_io_b = io_pp_17[4]; // @[wallaced.scala 89:18]
  assign FullAdder_122_io_ci = io_pp_18[3]; // @[wallaced.scala 90:19]
  assign FullAdder_123_io_a = io_pp_3[1]; // @[wallaced.scala 88:18]
  assign FullAdder_123_io_b = io_pp_4[0]; // @[wallaced.scala 89:18]
  assign FullAdder_123_io_ci = io_pp_16[4]; // @[wallaced.scala 90:19]
  assign FullAdder_124_io_a = io_pp_3[0]; // @[wallaced.scala 88:18]
  assign FullAdder_124_io_b = io_pp_16[3]; // @[wallaced.scala 89:18]
  assign FullAdder_124_io_ci = io_pp_17[2]; // @[wallaced.scala 90:19]
  assign FullAdder_125_io_a = io_pp_29[15]; // @[wallaced.scala 88:18]
  assign FullAdder_125_io_b = io_pp_30[14]; // @[wallaced.scala 89:18]
  assign FullAdder_125_io_ci = io_pp_31[13]; // @[wallaced.scala 90:19]
  assign FullAdder_126_io_a = io_pp_28[14]; // @[wallaced.scala 88:18]
  assign FullAdder_126_io_b = io_pp_29[13]; // @[wallaced.scala 89:18]
  assign FullAdder_126_io_ci = io_pp_30[12]; // @[wallaced.scala 90:19]
  assign FullAdder_127_io_a = io_pp_29[12]; // @[wallaced.scala 88:18]
  assign FullAdder_127_io_b = io_pp_30[11]; // @[wallaced.scala 89:18]
  assign FullAdder_127_io_ci = io_pp_31[10]; // @[wallaced.scala 90:19]
  assign FullAdder_128_io_a = io_pp_27[13]; // @[wallaced.scala 88:18]
  assign FullAdder_128_io_b = io_pp_28[12]; // @[wallaced.scala 89:18]
  assign FullAdder_128_io_ci = io_pp_29[11]; // @[wallaced.scala 90:19]
  assign FullAdder_129_io_a = io_pp_28[11]; // @[wallaced.scala 88:18]
  assign FullAdder_129_io_b = io_pp_29[10]; // @[wallaced.scala 89:18]
  assign FullAdder_129_io_ci = io_pp_30[9]; // @[wallaced.scala 90:19]
  assign FullAdder_130_io_a = io_pp_29[9]; // @[wallaced.scala 88:18]
  assign FullAdder_130_io_b = io_pp_30[8]; // @[wallaced.scala 89:18]
  assign FullAdder_130_io_ci = io_pp_31[7]; // @[wallaced.scala 90:19]
  assign FullAdder_131_io_a = io_pp_27[10]; // @[wallaced.scala 88:18]
  assign FullAdder_131_io_b = io_pp_28[9]; // @[wallaced.scala 89:18]
  assign FullAdder_131_io_ci = io_pp_29[8]; // @[wallaced.scala 90:19]
  assign FullAdder_132_io_a = io_pp_30[7]; // @[wallaced.scala 88:18]
  assign FullAdder_132_io_b = io_pp_31[6]; // @[wallaced.scala 89:18]
  assign FullAdder_132_io_ci = FullAdder_12_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_133_io_a = io_pp_28[8]; // @[wallaced.scala 88:18]
  assign FullAdder_133_io_b = io_pp_29[7]; // @[wallaced.scala 89:18]
  assign FullAdder_133_io_ci = io_pp_30[6]; // @[wallaced.scala 90:19]
  assign FullAdder_134_io_a = io_pp_26[9]; // @[wallaced.scala 88:18]
  assign FullAdder_134_io_b = io_pp_27[8]; // @[wallaced.scala 89:18]
  assign FullAdder_134_io_ci = io_pp_28[7]; // @[wallaced.scala 90:19]
  assign FullAdder_135_io_a = io_pp_29[6]; // @[wallaced.scala 88:18]
  assign FullAdder_135_io_b = io_pp_30[5]; // @[wallaced.scala 89:18]
  assign FullAdder_135_io_ci = io_pp_31[4]; // @[wallaced.scala 90:19]
  assign FullAdder_136_io_a = io_pp_27[7]; // @[wallaced.scala 88:18]
  assign FullAdder_136_io_b = io_pp_28[6]; // @[wallaced.scala 89:18]
  assign FullAdder_136_io_ci = io_pp_29[5]; // @[wallaced.scala 90:19]
  assign FullAdder_137_io_a = io_pp_30[4]; // @[wallaced.scala 88:18]
  assign FullAdder_137_io_b = io_pp_31[3]; // @[wallaced.scala 89:18]
  assign FullAdder_137_io_ci = FullAdder_22_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_138_io_a = io_pp_25[8]; // @[wallaced.scala 88:18]
  assign FullAdder_138_io_b = io_pp_26[7]; // @[wallaced.scala 89:18]
  assign FullAdder_138_io_ci = io_pp_27[6]; // @[wallaced.scala 90:19]
  assign FullAdder_139_io_a = io_pp_28[5]; // @[wallaced.scala 88:18]
  assign FullAdder_139_io_b = io_pp_29[4]; // @[wallaced.scala 89:18]
  assign FullAdder_139_io_ci = io_pp_30[3]; // @[wallaced.scala 90:19]
  assign FullAdder_140_io_a = io_pp_26[6]; // @[wallaced.scala 88:18]
  assign FullAdder_140_io_b = io_pp_27[5]; // @[wallaced.scala 89:18]
  assign FullAdder_140_io_ci = io_pp_28[4]; // @[wallaced.scala 90:19]
  assign FullAdder_141_io_a = io_pp_29[3]; // @[wallaced.scala 88:18]
  assign FullAdder_141_io_b = io_pp_30[2]; // @[wallaced.scala 89:18]
  assign FullAdder_141_io_ci = io_pp_31[1]; // @[wallaced.scala 90:19]
  assign FullAdder_142_io_a = io_pp_24[7]; // @[wallaced.scala 88:18]
  assign FullAdder_142_io_b = io_pp_25[6]; // @[wallaced.scala 89:18]
  assign FullAdder_142_io_ci = io_pp_26[5]; // @[wallaced.scala 90:19]
  assign FullAdder_143_io_a = io_pp_27[4]; // @[wallaced.scala 88:18]
  assign FullAdder_143_io_b = io_pp_28[3]; // @[wallaced.scala 89:18]
  assign FullAdder_143_io_ci = io_pp_29[2]; // @[wallaced.scala 90:19]
  assign FullAdder_144_io_a = io_pp_25[5]; // @[wallaced.scala 88:18]
  assign FullAdder_144_io_b = io_pp_26[4]; // @[wallaced.scala 89:18]
  assign FullAdder_144_io_ci = io_pp_27[3]; // @[wallaced.scala 90:19]
  assign FullAdder_145_io_a = io_pp_28[2]; // @[wallaced.scala 88:18]
  assign FullAdder_145_io_b = io_pp_29[1]; // @[wallaced.scala 89:18]
  assign FullAdder_145_io_ci = io_pp_30[0]; // @[wallaced.scala 90:19]
  assign FullAdder_146_io_a = io_pp_23[6]; // @[wallaced.scala 88:18]
  assign FullAdder_146_io_b = io_pp_24[5]; // @[wallaced.scala 89:18]
  assign FullAdder_146_io_ci = io_pp_25[4]; // @[wallaced.scala 90:19]
  assign FullAdder_147_io_a = io_pp_26[3]; // @[wallaced.scala 88:18]
  assign FullAdder_147_io_b = io_pp_27[2]; // @[wallaced.scala 89:18]
  assign FullAdder_147_io_ci = io_pp_28[1]; // @[wallaced.scala 90:19]
  assign FullAdder_148_io_a = io_pp_24[4]; // @[wallaced.scala 88:18]
  assign FullAdder_148_io_b = io_pp_25[3]; // @[wallaced.scala 89:18]
  assign FullAdder_148_io_ci = io_pp_26[2]; // @[wallaced.scala 90:19]
  assign FullAdder_149_io_a = io_pp_22[5]; // @[wallaced.scala 88:18]
  assign FullAdder_149_io_b = io_pp_23[4]; // @[wallaced.scala 89:18]
  assign FullAdder_149_io_ci = io_pp_24[3]; // @[wallaced.scala 90:19]
  assign FullAdder_150_io_a = io_pp_20[6]; // @[wallaced.scala 88:18]
  assign FullAdder_150_io_b = io_pp_21[5]; // @[wallaced.scala 89:18]
  assign FullAdder_150_io_ci = io_pp_22[4]; // @[wallaced.scala 90:19]
  assign FullAdder_151_io_a = io_pp_23[3]; // @[wallaced.scala 88:18]
  assign FullAdder_151_io_b = io_pp_24[2]; // @[wallaced.scala 89:18]
  assign FullAdder_151_io_ci = io_pp_25[1]; // @[wallaced.scala 90:19]
  assign FullAdder_152_io_a = io_pp_21[4]; // @[wallaced.scala 88:18]
  assign FullAdder_152_io_b = io_pp_22[3]; // @[wallaced.scala 89:18]
  assign FullAdder_152_io_ci = io_pp_23[2]; // @[wallaced.scala 90:19]
  assign FullAdder_153_io_a = io_pp_19[5]; // @[wallaced.scala 88:18]
  assign FullAdder_153_io_b = io_pp_20[4]; // @[wallaced.scala 89:18]
  assign FullAdder_153_io_ci = io_pp_21[3]; // @[wallaced.scala 90:19]
  assign HalfAdder_io_a = io_pp_22[2]; // @[wallaced.scala 79:18]
  assign HalfAdder_io_b = io_pp_23[1]; // @[wallaced.scala 80:18]
  assign FullAdder_154_io_a = io_pp_20[3]; // @[wallaced.scala 88:18]
  assign FullAdder_154_io_b = io_pp_21[2]; // @[wallaced.scala 89:18]
  assign FullAdder_154_io_ci = io_pp_22[1]; // @[wallaced.scala 90:19]
  assign FullAdder_155_io_a = io_pp_18[4]; // @[wallaced.scala 88:18]
  assign FullAdder_155_io_b = io_pp_19[3]; // @[wallaced.scala 89:18]
  assign FullAdder_155_io_ci = io_pp_20[2]; // @[wallaced.scala 90:19]
  assign FullAdder_156_io_a = io_pp_17[3]; // @[wallaced.scala 88:18]
  assign FullAdder_156_io_b = io_pp_18[2]; // @[wallaced.scala 89:18]
  assign FullAdder_156_io_ci = io_pp_19[1]; // @[wallaced.scala 90:19]
  assign FullAdder_157_io_a = io_pp_30[13]; // @[wallaced.scala 88:18]
  assign FullAdder_157_io_b = io_pp_31[12]; // @[wallaced.scala 89:18]
  assign FullAdder_157_io_ci = FullAdder_1_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_158_io_a = io_pp_31[11]; // @[wallaced.scala 88:18]
  assign FullAdder_158_io_b = FullAdder_2_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_158_io_ci = FullAdder_3_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_159_io_a = io_pp_30[10]; // @[wallaced.scala 88:18]
  assign FullAdder_159_io_b = io_pp_31[9]; // @[wallaced.scala 89:18]
  assign FullAdder_159_io_ci = FullAdder_5_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_160_io_a = io_pp_31[8]; // @[wallaced.scala 88:18]
  assign FullAdder_160_io_b = FullAdder_7_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_160_io_ci = FullAdder_8_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_161_io_a = FullAdder_9_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_161_io_b = FullAdder_10_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_161_io_ci = FullAdder_11_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_162_io_a = FullAdder_13_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_162_io_b = FullAdder_14_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_162_io_ci = FullAdder_15_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_163_io_a = io_pp_31[5]; // @[wallaced.scala 88:18]
  assign FullAdder_163_io_b = FullAdder_15_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_163_io_ci = FullAdder_16_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_164_io_a = FullAdder_18_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_164_io_b = FullAdder_19_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_164_io_ci = FullAdder_20_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_165_io_a = FullAdder_23_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_165_io_b = FullAdder_24_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_165_io_ci = FullAdder_25_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_166_io_a = io_pp_31[2]; // @[wallaced.scala 88:18]
  assign FullAdder_166_io_b = FullAdder_26_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_166_io_ci = FullAdder_27_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_167_io_a = FullAdder_28_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_167_io_b = FullAdder_29_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_167_io_ci = FullAdder_30_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_168_io_a = FullAdder_30_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_168_io_b = FullAdder_31_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_168_io_ci = FullAdder_32_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_169_io_a = io_pp_30[1]; // @[wallaced.scala 88:18]
  assign FullAdder_169_io_b = io_pp_31[0]; // @[wallaced.scala 89:18]
  assign FullAdder_169_io_ci = FullAdder_35_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_170_io_a = FullAdder_36_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_170_io_b = FullAdder_37_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_170_io_ci = FullAdder_38_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_171_io_a = FullAdder_40_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_171_io_b = FullAdder_41_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_171_io_ci = FullAdder_42_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_172_io_a = io_pp_29[0]; // @[wallaced.scala 88:18]
  assign FullAdder_172_io_b = FullAdder_45_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_172_io_ci = FullAdder_46_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_173_io_a = io_pp_27[1]; // @[wallaced.scala 88:18]
  assign FullAdder_173_io_b = io_pp_28[0]; // @[wallaced.scala 89:18]
  assign FullAdder_173_io_ci = FullAdder_49_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_174_io_a = io_pp_25[2]; // @[wallaced.scala 88:18]
  assign FullAdder_174_io_b = io_pp_26[1]; // @[wallaced.scala 89:18]
  assign FullAdder_174_io_ci = io_pp_27[0]; // @[wallaced.scala 90:19]
  assign HalfAdder_1_io_a = FullAdder_53_io_s; // @[wallaced.scala 79:18]
  assign HalfAdder_1_io_b = FullAdder_54_io_s; // @[wallaced.scala 80:18]
  assign FullAdder_175_io_a = io_pp_26[0]; // @[wallaced.scala 88:18]
  assign FullAdder_175_io_b = FullAdder_57_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_175_io_ci = FullAdder_58_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_176_io_a = io_pp_24[1]; // @[wallaced.scala 88:18]
  assign FullAdder_176_io_b = io_pp_25[0]; // @[wallaced.scala 89:18]
  assign FullAdder_176_io_ci = FullAdder_60_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_177_io_a = io_pp_24[0]; // @[wallaced.scala 88:18]
  assign FullAdder_177_io_b = FullAdder_63_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_177_io_ci = FullAdder_64_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_178_io_a = io_pp_19[2]; // @[wallaced.scala 88:18]
  assign FullAdder_178_io_b = io_pp_20[1]; // @[wallaced.scala 89:18]
  assign FullAdder_178_io_ci = io_pp_21[0]; // @[wallaced.scala 90:19]
  assign FullAdder_179_io_a = FullAdder_3_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_179_io_b = FullAdder_4_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_179_io_ci = FullAdder_5_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_180_io_a = FullAdder_6_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_180_io_b = FullAdder_7_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_180_io_ci = FullAdder_8_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_181_io_a = FullAdder_9_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_181_io_b = FullAdder_10_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_181_io_ci = FullAdder_11_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_182_io_a = FullAdder_12_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_182_io_b = FullAdder_13_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_182_io_ci = FullAdder_14_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_183_io_a = FullAdder_17_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_183_io_b = FullAdder_18_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_183_io_ci = FullAdder_19_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_184_io_a = FullAdder_21_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_184_io_b = FullAdder_22_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_184_io_ci = FullAdder_23_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_185_io_a = FullAdder_26_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_185_io_b = FullAdder_27_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_185_io_ci = FullAdder_28_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_186_io_a = FullAdder_31_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_186_io_b = FullAdder_32_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_186_io_ci = FullAdder_33_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_187_io_a = FullAdder_33_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_187_io_b = FullAdder_34_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_187_io_ci = FullAdder_35_io_co; // @[wallaced.scala 90:19]
  assign HalfAdder_2_io_a = FullAdder_36_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_2_io_b = FullAdder_37_io_co; // @[wallaced.scala 80:18]
  assign FullAdder_188_io_a = FullAdder_39_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_188_io_b = FullAdder_40_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_188_io_ci = FullAdder_41_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_189_io_a = FullAdder_43_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_189_io_b = FullAdder_44_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_189_io_ci = FullAdder_45_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_190_io_a = FullAdder_47_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_190_io_b = FullAdder_48_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_190_io_ci = FullAdder_49_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_191_io_a = FullAdder_50_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_191_io_b = FullAdder_51_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_191_io_ci = FullAdder_52_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_192_io_a = FullAdder_55_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_192_io_b = FullAdder_56_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_192_io_ci = FullAdder_57_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_193_io_a = FullAdder_61_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_193_io_b = FullAdder_62_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_193_io_ci = FullAdder_63_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_194_io_a = io_pp_21[1]; // @[wallaced.scala 88:18]
  assign FullAdder_194_io_b = io_pp_22[0]; // @[wallaced.scala 89:18]
  assign FullAdder_194_io_ci = FullAdder_68_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_195_io_a = FullAdder_16_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_195_io_b = FullAdder_17_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_195_io_ci = FullAdder_84_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_196_io_a = FullAdder_20_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_196_io_b = FullAdder_21_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_196_io_ci = FullAdder_86_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_197_io_a = FullAdder_24_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_197_io_b = FullAdder_25_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_197_io_ci = FullAdder_89_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_198_io_a = FullAdder_29_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_198_io_b = FullAdder_91_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_198_io_ci = FullAdder_92_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_199_io_a = FullAdder_34_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_199_io_b = FullAdder_94_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_199_io_ci = FullAdder_95_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_200_io_a = FullAdder_38_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_200_io_b = FullAdder_39_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_200_io_ci = FullAdder_97_io_s; // @[wallaced.scala 90:19]
  assign HalfAdder_3_io_a = FullAdder_42_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_3_io_b = FullAdder_43_io_co; // @[wallaced.scala 80:18]
  assign HalfAdder_4_io_a = FullAdder_46_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_4_io_b = FullAdder_47_io_co; // @[wallaced.scala 80:18]
  assign HalfAdder_5_io_a = FullAdder_50_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_5_io_b = FullAdder_51_io_co; // @[wallaced.scala 80:18]
  assign FullAdder_201_io_a = FullAdder_53_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_201_io_b = FullAdder_54_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_201_io_ci = FullAdder_55_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_202_io_a = FullAdder_59_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_202_io_b = FullAdder_60_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_202_io_ci = FullAdder_61_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_203_io_a = io_pp_23[0]; // @[wallaced.scala 88:18]
  assign FullAdder_203_io_b = FullAdder_66_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_203_io_ci = FullAdder_67_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_204_io_a = FullAdder_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_204_io_b = FullAdder_1_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_204_io_ci = FullAdder_76_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_205_io_a = FullAdder_2_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_205_io_b = FullAdder_76_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_205_io_ci = FullAdder_77_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_206_io_a = FullAdder_4_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_206_io_b = FullAdder_77_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_206_io_ci = FullAdder_78_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_207_io_a = FullAdder_6_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_207_io_b = FullAdder_78_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_207_io_ci = FullAdder_79_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_208_io_a = FullAdder_127_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_208_io_b = FullAdder_128_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_208_io_ci = FullAdder_159_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_209_io_a = FullAdder_79_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_209_io_b = FullAdder_80_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_209_io_ci = FullAdder_81_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_210_io_a = FullAdder_128_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_210_io_b = FullAdder_129_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_210_io_ci = FullAdder_159_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_211_io_a = FullAdder_80_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_211_io_b = FullAdder_81_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_211_io_ci = FullAdder_82_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_212_io_a = FullAdder_83_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_212_io_b = FullAdder_129_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_212_io_ci = FullAdder_130_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_213_io_a = FullAdder_82_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_213_io_b = FullAdder_83_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_213_io_ci = FullAdder_84_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_214_io_a = FullAdder_85_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_214_io_b = FullAdder_130_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_214_io_ci = FullAdder_131_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_215_io_a = FullAdder_132_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_215_io_b = FullAdder_161_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_215_io_ci = FullAdder_162_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_216_io_a = FullAdder_85_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_216_io_b = FullAdder_86_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_216_io_ci = FullAdder_87_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_217_io_a = FullAdder_88_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_217_io_b = FullAdder_131_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_217_io_ci = FullAdder_132_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_218_io_a = FullAdder_133_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_218_io_b = FullAdder_162_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_218_io_ci = FullAdder_163_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_219_io_a = FullAdder_87_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_219_io_b = FullAdder_88_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_219_io_ci = FullAdder_89_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_220_io_a = FullAdder_90_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_220_io_b = FullAdder_133_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_220_io_ci = FullAdder_134_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_221_io_a = FullAdder_135_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_221_io_b = FullAdder_163_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_221_io_ci = FullAdder_164_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_222_io_a = FullAdder_90_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_222_io_b = FullAdder_91_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_222_io_ci = FullAdder_92_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_223_io_a = FullAdder_93_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_223_io_b = FullAdder_134_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_223_io_ci = FullAdder_135_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_224_io_a = FullAdder_136_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_224_io_b = FullAdder_137_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_224_io_ci = FullAdder_164_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_225_io_a = FullAdder_165_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_225_io_b = FullAdder_184_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_225_io_ci = FullAdder_185_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_226_io_a = FullAdder_93_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_226_io_b = FullAdder_94_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_226_io_ci = FullAdder_95_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_227_io_a = FullAdder_96_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_227_io_b = FullAdder_136_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_227_io_ci = FullAdder_137_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_228_io_a = FullAdder_138_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_228_io_b = FullAdder_139_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_228_io_ci = FullAdder_165_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_229_io_a = FullAdder_166_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_229_io_b = FullAdder_167_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_229_io_ci = FullAdder_185_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_230_io_a = FullAdder_96_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_230_io_b = FullAdder_97_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_230_io_ci = FullAdder_98_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_231_io_a = FullAdder_99_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_231_io_b = FullAdder_138_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_231_io_ci = FullAdder_139_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_232_io_a = FullAdder_140_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_232_io_b = FullAdder_141_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_232_io_ci = FullAdder_166_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_233_io_a = FullAdder_167_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_233_io_b = FullAdder_168_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_233_io_ci = FullAdder_186_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_234_io_a = FullAdder_98_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_234_io_b = FullAdder_99_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_234_io_ci = FullAdder_100_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_235_io_a = FullAdder_101_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_235_io_b = FullAdder_102_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_235_io_ci = FullAdder_140_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_236_io_a = FullAdder_141_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_236_io_b = FullAdder_142_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_236_io_ci = FullAdder_143_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_237_io_a = FullAdder_168_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_237_io_b = FullAdder_169_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_237_io_ci = FullAdder_170_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_238_io_a = FullAdder_187_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_238_io_b = HalfAdder_2_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_238_io_ci = FullAdder_188_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_239_io_a = FullAdder_44_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_239_io_b = FullAdder_100_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_239_io_ci = FullAdder_101_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_240_io_a = FullAdder_102_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_240_io_b = FullAdder_103_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_240_io_ci = FullAdder_104_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_241_io_a = FullAdder_105_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_241_io_b = FullAdder_142_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_241_io_ci = FullAdder_143_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_242_io_a = FullAdder_144_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_242_io_b = FullAdder_145_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_242_io_ci = FullAdder_169_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_243_io_a = FullAdder_170_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_243_io_b = FullAdder_171_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_243_io_ci = FullAdder_188_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_244_io_a = FullAdder_48_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_244_io_b = FullAdder_103_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_244_io_ci = FullAdder_104_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_245_io_a = FullAdder_105_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_245_io_b = FullAdder_106_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_245_io_ci = FullAdder_107_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_246_io_a = FullAdder_108_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_246_io_b = FullAdder_144_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_246_io_ci = FullAdder_145_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_247_io_a = FullAdder_146_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_247_io_b = FullAdder_147_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_247_io_ci = FullAdder_171_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_248_io_a = FullAdder_172_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_248_io_b = FullAdder_189_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_248_io_ci = FullAdder_190_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_249_io_a = FullAdder_52_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_249_io_b = FullAdder_106_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_249_io_ci = FullAdder_107_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_250_io_a = FullAdder_108_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_250_io_b = FullAdder_109_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_250_io_ci = FullAdder_110_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_251_io_a = FullAdder_111_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_251_io_b = FullAdder_146_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_251_io_ci = FullAdder_147_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_252_io_a = FullAdder_148_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_252_io_b = FullAdder_172_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_252_io_ci = FullAdder_173_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_253_io_a = FullAdder_56_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_253_io_b = FullAdder_109_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_253_io_ci = FullAdder_110_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_254_io_a = FullAdder_111_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_254_io_b = FullAdder_112_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_254_io_ci = FullAdder_113_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_255_io_a = FullAdder_148_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_255_io_b = FullAdder_149_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_255_io_ci = FullAdder_173_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_256_io_a = FullAdder_174_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_256_io_b = HalfAdder_1_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_256_io_ci = FullAdder_191_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_257_io_a = FullAdder_58_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_257_io_b = FullAdder_59_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_257_io_ci = FullAdder_112_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_258_io_a = FullAdder_113_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_258_io_b = FullAdder_114_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_258_io_ci = FullAdder_115_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_259_io_a = FullAdder_149_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_259_io_b = FullAdder_150_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_259_io_ci = FullAdder_151_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_260_io_a = FullAdder_174_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_260_io_b = HalfAdder_1_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_260_io_ci = FullAdder_175_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_261_io_a = FullAdder_62_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_261_io_b = FullAdder_114_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_261_io_ci = FullAdder_115_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_262_io_a = FullAdder_116_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_262_io_b = FullAdder_117_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_262_io_ci = FullAdder_150_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_263_io_a = FullAdder_151_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_263_io_b = FullAdder_152_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_263_io_ci = FullAdder_175_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_264_io_a = FullAdder_64_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_264_io_b = FullAdder_65_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_264_io_ci = FullAdder_116_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_265_io_a = FullAdder_117_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_265_io_b = FullAdder_118_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_265_io_ci = FullAdder_152_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_266_io_a = FullAdder_153_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_266_io_b = HalfAdder_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_266_io_ci = FullAdder_176_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_267_io_a = FullAdder_65_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_267_io_b = FullAdder_66_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_267_io_ci = FullAdder_67_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_268_io_a = FullAdder_118_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_268_io_b = FullAdder_119_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_268_io_ci = FullAdder_120_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_269_io_a = FullAdder_153_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_269_io_b = HalfAdder_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_269_io_ci = FullAdder_154_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_270_io_a = FullAdder_68_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_270_io_b = FullAdder_69_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_270_io_ci = FullAdder_119_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_271_io_a = FullAdder_120_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_271_io_b = FullAdder_121_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_271_io_ci = FullAdder_154_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_272_io_a = FullAdder_69_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_272_io_b = FullAdder_70_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_272_io_ci = FullAdder_71_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_273_io_a = FullAdder_121_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_273_io_b = FullAdder_122_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_273_io_ci = FullAdder_155_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_274_io_a = FullAdder_70_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_274_io_b = FullAdder_71_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_274_io_ci = FullAdder_72_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_275_io_a = FullAdder_122_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_275_io_b = FullAdder_123_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_275_io_ci = FullAdder_156_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_276_io_a = io_pp_20[0]; // @[wallaced.scala 88:18]
  assign FullAdder_276_io_b = FullAdder_72_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_276_io_ci = FullAdder_73_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_277_io_a = io_pp_18[1]; // @[wallaced.scala 88:18]
  assign FullAdder_277_io_b = io_pp_19[0]; // @[wallaced.scala 89:18]
  assign FullAdder_277_io_ci = FullAdder_73_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_278_io_a = io_pp_16[2]; // @[wallaced.scala 88:18]
  assign FullAdder_278_io_b = io_pp_17[1]; // @[wallaced.scala 89:18]
  assign FullAdder_278_io_ci = io_pp_18[0]; // @[wallaced.scala 90:19]
  assign FullAdder_279_io_a = io_pp_31[14]; // @[wallaced.scala 88:18]
  assign FullAdder_279_io_b = FullAdder_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_279_io_ci = FullAdder_75_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_280_io_a = FullAdder_126_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_280_io_b = FullAdder_157_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_280_io_ci = FullAdder_158_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_281_io_a = FullAdder_126_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_281_io_b = FullAdder_127_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_281_io_ci = FullAdder_158_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_282_io_a = FullAdder_179_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_282_io_b = FullAdder_180_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_282_io_ci = FullAdder_207_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_283_io_a = FullAdder_160_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_283_io_b = FullAdder_180_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_283_io_ci = FullAdder_181_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_284_io_a = FullAdder_160_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_284_io_b = FullAdder_161_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_284_io_ci = FullAdder_181_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_285_io_a = FullAdder_182_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_285_io_b = FullAdder_211_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_285_io_ci = FullAdder_212_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_286_io_a = FullAdder_182_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_286_io_b = FullAdder_195_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_286_io_ci = FullAdder_213_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_287_io_a = FullAdder_214_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_287_io_b = FullAdder_215_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_287_io_ci = FullAdder_216_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_288_io_a = FullAdder_183_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_288_io_b = FullAdder_195_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_288_io_ci = FullAdder_196_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_289_io_a = FullAdder_216_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_289_io_b = FullAdder_217_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_289_io_ci = FullAdder_218_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_290_io_a = FullAdder_183_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_290_io_b = FullAdder_184_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_290_io_ci = FullAdder_196_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_291_io_a = FullAdder_197_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_291_io_b = FullAdder_219_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_291_io_ci = FullAdder_220_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_292_io_a = FullAdder_221_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_292_io_b = FullAdder_222_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_292_io_ci = FullAdder_223_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_293_io_a = FullAdder_197_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_293_io_b = FullAdder_198_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_293_io_ci = FullAdder_222_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_294_io_a = FullAdder_223_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_294_io_b = FullAdder_224_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_294_io_ci = FullAdder_225_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_295_io_a = FullAdder_186_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_295_io_b = FullAdder_198_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_295_io_ci = FullAdder_199_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_296_io_a = FullAdder_226_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_296_io_b = FullAdder_227_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_296_io_ci = FullAdder_228_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_297_io_a = FullAdder_229_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_297_io_b = FullAdder_230_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_297_io_ci = FullAdder_231_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_298_io_a = FullAdder_187_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_298_io_b = HalfAdder_2_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_298_io_ci = FullAdder_199_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_299_io_a = FullAdder_200_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_299_io_b = FullAdder_230_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_299_io_ci = FullAdder_231_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_300_io_a = FullAdder_232_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_300_io_b = FullAdder_233_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_300_io_ci = FullAdder_234_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_301_io_a = FullAdder_200_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_301_io_b = HalfAdder_3_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_301_io_ci = FullAdder_234_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_302_io_a = FullAdder_235_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_302_io_b = FullAdder_236_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_302_io_ci = FullAdder_237_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_303_io_a = FullAdder_238_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_303_io_b = FullAdder_239_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_303_io_ci = FullAdder_240_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_304_io_a = FullAdder_189_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_304_io_b = HalfAdder_3_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_304_io_ci = HalfAdder_4_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_305_io_a = FullAdder_239_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_305_io_b = FullAdder_240_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_305_io_ci = FullAdder_241_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_306_io_a = FullAdder_242_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_306_io_b = FullAdder_243_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_306_io_ci = FullAdder_244_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_307_io_a = HalfAdder_4_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_307_io_b = HalfAdder_5_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_307_io_ci = FullAdder_244_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_308_io_a = FullAdder_245_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_308_io_b = FullAdder_246_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_308_io_ci = FullAdder_247_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_309_io_a = FullAdder_248_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_309_io_b = FullAdder_249_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_309_io_ci = FullAdder_250_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_310_io_a = FullAdder_190_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_310_io_b = FullAdder_191_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_310_io_ci = HalfAdder_5_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_311_io_a = FullAdder_201_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_311_io_b = FullAdder_249_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_311_io_ci = FullAdder_250_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_312_io_a = FullAdder_251_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_312_io_b = FullAdder_252_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_312_io_ci = FullAdder_253_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_313_io_a = FullAdder_192_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_313_io_b = FullAdder_201_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_313_io_ci = FullAdder_253_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_314_io_a = FullAdder_254_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_314_io_b = FullAdder_255_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_314_io_ci = FullAdder_256_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_315_io_a = FullAdder_257_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_315_io_b = FullAdder_258_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_315_io_ci = FullAdder_259_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_316_io_a = FullAdder_192_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_316_io_b = FullAdder_202_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_316_io_ci = FullAdder_257_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_317_io_a = FullAdder_258_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_317_io_b = FullAdder_259_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_317_io_ci = FullAdder_260_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_318_io_a = FullAdder_176_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_318_io_b = FullAdder_193_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_318_io_ci = FullAdder_202_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_319_io_a = FullAdder_261_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_319_io_b = FullAdder_262_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_319_io_ci = FullAdder_263_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_320_io_a = FullAdder_177_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_320_io_b = FullAdder_193_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_320_io_ci = FullAdder_264_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_321_io_a = FullAdder_265_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_321_io_b = FullAdder_266_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_321_io_ci = FullAdder_267_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_322_io_a = FullAdder_177_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_322_io_b = FullAdder_203_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_322_io_ci = FullAdder_267_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_323_io_a = FullAdder_155_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_323_io_b = FullAdder_194_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_323_io_ci = FullAdder_203_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_324_io_a = FullAdder_270_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_324_io_b = FullAdder_271_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_324_io_ci = FullAdder_272_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_325_io_a = FullAdder_178_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_325_io_b = FullAdder_194_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_325_io_ci = FullAdder_272_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_326_io_a = FullAdder_178_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_326_io_b = FullAdder_274_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_326_io_ci = FullAdder_275_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_327_io_a = FullAdder_123_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_327_io_b = FullAdder_124_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_327_io_ci = FullAdder_156_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_328_io_a = FullAdder_74_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_328_io_b = FullAdder_124_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_328_io_ci = FullAdder_277_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_329_io_a = FullAdder_125_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_329_io_b = FullAdder_157_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_329_io_ci = FullAdder_204_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_330_io_a = FullAdder_179_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_330_io_b = FullAdder_206_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_330_io_ci = FullAdder_207_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_331_io_a = FullAdder_208_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_331_io_b = FullAdder_209_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_331_io_ci = FullAdder_210_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_332_io_a = FullAdder_209_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_332_io_b = FullAdder_210_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_332_io_ci = FullAdder_211_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_333_io_a = FullAdder_213_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_333_io_b = FullAdder_214_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_333_io_ci = FullAdder_215_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_334_io_a = FullAdder_217_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_334_io_b = FullAdder_218_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_334_io_ci = FullAdder_286_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_335_io_a = FullAdder_219_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_335_io_b = FullAdder_220_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_335_io_ci = FullAdder_221_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_336_io_a = FullAdder_288_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_336_io_b = FullAdder_289_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_336_io_ci = FullAdder_290_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_337_io_a = FullAdder_224_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_337_io_b = FullAdder_225_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_337_io_ci = FullAdder_290_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_338_io_a = FullAdder_226_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_338_io_b = FullAdder_227_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_338_io_ci = FullAdder_228_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_339_io_a = FullAdder_229_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_339_io_b = FullAdder_293_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_339_io_ci = FullAdder_294_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_340_io_a = FullAdder_232_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_340_io_b = FullAdder_233_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_340_io_ci = FullAdder_295_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_341_io_a = FullAdder_296_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_341_io_b = FullAdder_297_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_341_io_ci = FullAdder_298_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_342_io_a = FullAdder_235_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_342_io_b = FullAdder_236_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_342_io_ci = FullAdder_237_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_343_io_a = FullAdder_238_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_343_io_b = FullAdder_298_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_343_io_ci = FullAdder_299_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_344_io_a = FullAdder_241_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_344_io_b = FullAdder_242_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_344_io_ci = FullAdder_243_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_345_io_a = FullAdder_301_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_345_io_b = FullAdder_302_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_345_io_ci = FullAdder_303_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_346_io_a = FullAdder_245_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_346_io_b = FullAdder_246_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_346_io_ci = FullAdder_247_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_347_io_a = FullAdder_248_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_347_io_b = FullAdder_304_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_347_io_ci = FullAdder_305_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_348_io_a = FullAdder_251_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_348_io_b = FullAdder_252_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_348_io_ci = FullAdder_307_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_349_io_a = FullAdder_308_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_349_io_b = FullAdder_309_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_349_io_ci = FullAdder_310_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_350_io_a = FullAdder_254_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_350_io_b = FullAdder_255_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_350_io_ci = FullAdder_256_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_351_io_a = FullAdder_310_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_351_io_b = FullAdder_311_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_351_io_ci = FullAdder_312_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_352_io_a = FullAdder_260_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_352_io_b = FullAdder_313_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_352_io_ci = FullAdder_314_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_353_io_a = FullAdder_261_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_353_io_b = FullAdder_262_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_353_io_ci = FullAdder_263_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_354_io_a = FullAdder_264_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_354_io_b = FullAdder_265_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_354_io_ci = FullAdder_266_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_355_io_a = FullAdder_318_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_355_io_b = FullAdder_319_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_355_io_ci = FullAdder_320_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_356_io_a = FullAdder_268_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_356_io_b = FullAdder_269_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_356_io_ci = FullAdder_320_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_357_io_a = FullAdder_268_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_357_io_b = FullAdder_269_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_357_io_ci = FullAdder_270_io_co; // @[wallaced.scala 90:19]
  assign HalfAdder_6_io_a = FullAdder_271_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_6_io_b = FullAdder_322_io_s; // @[wallaced.scala 80:18]
  assign FullAdder_358_io_a = FullAdder_273_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_358_io_b = FullAdder_323_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_358_io_ci = FullAdder_324_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_359_io_a = FullAdder_273_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_359_io_b = FullAdder_274_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_359_io_ci = FullAdder_275_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_360_io_a = FullAdder_276_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_360_io_b = FullAdder_277_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_360_io_ci = FullAdder_327_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_361_io_a = FullAdder_205_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_361_io_b = FullAdder_206_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_361_io_ci = FullAdder_280_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_362_io_a = FullAdder_208_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_362_io_b = FullAdder_281_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_362_io_ci = FullAdder_282_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_363_io_a = FullAdder_212_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_363_io_b = FullAdder_283_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_363_io_ci = FullAdder_284_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_364_io_a = FullAdder_284_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_364_io_b = FullAdder_285_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_364_io_ci = FullAdder_286_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_365_io_a = FullAdder_287_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_365_io_b = FullAdder_288_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_365_io_ci = FullAdder_289_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_366_io_a = FullAdder_291_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_366_io_b = FullAdder_292_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_366_io_ci = FullAdder_335_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_367_io_a = FullAdder_291_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_367_io_b = FullAdder_292_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_367_io_ci = FullAdder_293_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_368_io_a = FullAdder_295_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_368_io_b = FullAdder_296_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_368_io_ci = FullAdder_297_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_369_io_a = FullAdder_299_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_369_io_b = FullAdder_300_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_369_io_ci = FullAdder_340_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_370_io_a = FullAdder_300_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_370_io_b = FullAdder_301_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_370_io_ci = FullAdder_302_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_371_io_a = FullAdder_303_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_371_io_b = FullAdder_342_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_371_io_ci = FullAdder_343_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_372_io_a = FullAdder_304_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_372_io_b = FullAdder_305_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_372_io_ci = FullAdder_306_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_373_io_a = FullAdder_306_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_373_io_b = FullAdder_307_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_373_io_ci = FullAdder_308_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_374_io_a = FullAdder_309_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_374_io_b = FullAdder_346_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_374_io_ci = FullAdder_347_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_375_io_a = FullAdder_311_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_375_io_b = FullAdder_312_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_375_io_ci = FullAdder_348_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_376_io_a = FullAdder_313_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_376_io_b = FullAdder_314_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_376_io_ci = FullAdder_315_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_377_io_a = FullAdder_315_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_377_io_b = FullAdder_316_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_377_io_ci = FullAdder_317_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_378_io_a = FullAdder_316_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_378_io_b = FullAdder_317_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_378_io_ci = FullAdder_318_io_co; // @[wallaced.scala 90:19]
  assign HalfAdder_7_io_a = FullAdder_319_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_7_io_b = FullAdder_353_io_s; // @[wallaced.scala 80:18]
  assign FullAdder_379_io_a = FullAdder_321_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_379_io_b = FullAdder_354_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_379_io_ci = FullAdder_355_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_380_io_a = FullAdder_321_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_380_io_b = FullAdder_322_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_380_io_ci = FullAdder_356_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_381_io_a = FullAdder_323_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_381_io_b = FullAdder_324_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_381_io_ci = FullAdder_357_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_382_io_a = FullAdder_276_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_382_io_b = FullAdder_326_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_382_io_ci = FullAdder_327_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_383_io_a = FullAdder_282_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_383_io_b = FullAdder_283_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_383_io_ci = FullAdder_331_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_384_io_a = FullAdder_285_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_384_io_b = FullAdder_332_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_384_io_ci = FullAdder_333_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_385_io_a = FullAdder_287_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_385_io_b = FullAdder_333_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_385_io_ci = FullAdder_334_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_386_io_a = FullAdder_334_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_386_io_b = FullAdder_335_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_386_io_ci = FullAdder_336_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_387_io_a = FullAdder_294_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_387_io_b = FullAdder_337_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_387_io_ci = FullAdder_338_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_388_io_a = FullAdder_338_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_388_io_b = FullAdder_339_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_388_io_ci = FullAdder_340_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_389_io_a = FullAdder_341_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_389_io_b = FullAdder_342_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_389_io_ci = FullAdder_343_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_390_io_a = FullAdder_344_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_390_io_b = FullAdder_345_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_390_io_ci = FullAdder_370_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_391_io_a = FullAdder_344_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_391_io_b = FullAdder_345_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_391_io_ci = FullAdder_346_io_co; // @[wallaced.scala 90:19]
  assign HalfAdder_8_io_a = FullAdder_347_io_co; // @[wallaced.scala 79:18]
  assign HalfAdder_8_io_b = FullAdder_372_io_s; // @[wallaced.scala 80:18]
  assign FullAdder_392_io_a = FullAdder_348_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_392_io_b = FullAdder_349_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_392_io_ci = FullAdder_373_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_393_io_a = FullAdder_349_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_393_io_b = FullAdder_350_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_393_io_ci = FullAdder_351_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_394_io_a = FullAdder_350_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_394_io_b = FullAdder_351_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_394_io_ci = FullAdder_352_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_395_io_a = FullAdder_352_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_395_io_b = FullAdder_353_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_395_io_ci = FullAdder_377_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_396_io_a = FullAdder_354_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_396_io_b = FullAdder_355_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_396_io_ci = FullAdder_378_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_397_io_a = FullAdder_357_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_397_io_b = HalfAdder_6_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_397_io_ci = FullAdder_380_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_398_io_a = FullAdder_325_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_398_io_b = FullAdder_326_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_398_io_ci = FullAdder_359_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_399_io_a = FullAdder_336_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_399_io_b = FullAdder_337_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_399_io_ci = FullAdder_366_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_400_io_a = FullAdder_339_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_400_io_b = FullAdder_367_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_400_io_ci = FullAdder_368_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_401_io_a = FullAdder_341_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_401_io_b = FullAdder_368_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_401_io_ci = FullAdder_369_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_402_io_a = FullAdder_369_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_402_io_b = FullAdder_370_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_402_io_ci = FullAdder_371_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_403_io_a = FullAdder_371_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_403_io_b = FullAdder_372_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_403_io_ci = FullAdder_390_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_404_io_a = FullAdder_373_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_404_io_b = FullAdder_374_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_404_io_ci = FullAdder_391_io_s; // @[wallaced.scala 90:19]
  assign HalfAdder_9_io_a = FullAdder_374_io_s; // @[wallaced.scala 79:18]
  assign HalfAdder_9_io_b = FullAdder_375_io_co; // @[wallaced.scala 80:18]
  assign HalfAdder_10_io_a = FullAdder_375_io_s; // @[wallaced.scala 79:18]
  assign HalfAdder_10_io_b = FullAdder_376_io_co; // @[wallaced.scala 80:18]
  assign HalfAdder_11_io_a = FullAdder_376_io_s; // @[wallaced.scala 79:18]
  assign HalfAdder_11_io_b = FullAdder_377_io_co; // @[wallaced.scala 80:18]
  assign FullAdder_405_io_a = FullAdder_378_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_405_io_b = HalfAdder_7_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_405_io_ci = FullAdder_395_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_406_io_a = FullAdder_356_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_406_io_b = FullAdder_379_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_406_io_ci = FullAdder_380_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_407_io_a = FullAdder_325_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_407_io_b = FullAdder_358_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_407_io_ci = FullAdder_359_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_408_io_a = io_pp_15[15]; // @[wallaced.scala 88:18]
  assign FullAdder_408_io_b = io_pp_31[15]; // @[wallaced.scala 89:18]
  assign FullAdder_408_io_ci = FullAdder_75_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_409_io_a = FullAdder_125_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_409_io_b = FullAdder_204_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_409_io_ci = FullAdder_279_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_410_io_a = FullAdder_205_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_410_io_b = FullAdder_280_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_410_io_ci = FullAdder_329_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_411_io_a = FullAdder_281_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_411_io_b = FullAdder_330_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_411_io_ci = FullAdder_361_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_412_io_a = FullAdder_330_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_412_io_b = FullAdder_331_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_412_io_ci = FullAdder_362_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_413_io_a = FullAdder_332_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_413_io_b = FullAdder_363_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_413_io_ci = FullAdder_383_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_414_io_a = FullAdder_363_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_414_io_b = FullAdder_364_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_414_io_ci = FullAdder_384_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_415_io_a = FullAdder_364_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_415_io_b = FullAdder_365_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_415_io_ci = FullAdder_385_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_416_io_a = FullAdder_365_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_416_io_b = FullAdder_366_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_416_io_ci = FullAdder_386_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_417_io_a = FullAdder_367_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_417_io_b = FullAdder_387_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_417_io_ci = FullAdder_399_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_418_io_a = FullAdder_387_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_418_io_b = FullAdder_388_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_418_io_ci = FullAdder_400_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_419_io_a = FullAdder_388_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_419_io_b = FullAdder_389_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_419_io_ci = FullAdder_401_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_420_io_a = FullAdder_389_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_420_io_b = FullAdder_390_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_420_io_ci = FullAdder_402_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_421_io_a = FullAdder_391_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_421_io_b = HalfAdder_8_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_421_io_ci = FullAdder_403_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_422_io_a = HalfAdder_8_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_422_io_b = FullAdder_392_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_422_io_ci = FullAdder_404_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_423_io_a = FullAdder_392_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_423_io_b = FullAdder_393_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_423_io_ci = HalfAdder_9_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_424_io_a = FullAdder_393_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_424_io_b = FullAdder_394_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_424_io_ci = HalfAdder_10_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_425_io_a = FullAdder_394_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_425_io_b = FullAdder_395_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_425_io_ci = HalfAdder_11_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_426_io_a = HalfAdder_7_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_426_io_b = FullAdder_379_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_426_io_ci = FullAdder_396_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_427_io_a = HalfAdder_6_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_427_io_b = FullAdder_358_io_co; // @[wallaced.scala 89:18]
  assign FullAdder_427_io_ci = FullAdder_381_io_s; // @[wallaced.scala 90:19]
  assign FullAdder_428_io_a = io_pp_0[1]; // @[wallaced.scala 88:18]
  assign FullAdder_428_io_b = io_pp_1[0]; // @[wallaced.scala 89:18]
  assign FullAdder_428_io_ci = io_pp_16[1]; // @[wallaced.scala 90:19]
  assign FullAdder_429_io_a = FullAdder_279_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_429_io_b = FullAdder_408_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_429_io_ci = FullAdder_409_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_430_io_a = FullAdder_329_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_430_io_b = FullAdder_409_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_430_io_ci = FullAdder_410_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_431_io_a = FullAdder_361_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_431_io_b = FullAdder_410_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_431_io_ci = FullAdder_411_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_432_io_a = FullAdder_362_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_432_io_b = FullAdder_411_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_432_io_ci = FullAdder_412_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_433_io_a = FullAdder_383_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_433_io_b = FullAdder_412_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_433_io_ci = FullAdder_413_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_434_io_a = FullAdder_384_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_434_io_b = FullAdder_413_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_434_io_ci = FullAdder_414_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_435_io_a = FullAdder_385_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_435_io_b = FullAdder_414_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_435_io_ci = FullAdder_415_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_436_io_a = FullAdder_386_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_436_io_b = FullAdder_415_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_436_io_ci = FullAdder_416_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_437_io_a = FullAdder_399_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_437_io_b = FullAdder_416_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_437_io_ci = FullAdder_417_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_438_io_a = FullAdder_400_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_438_io_b = FullAdder_417_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_438_io_ci = FullAdder_418_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_439_io_a = FullAdder_401_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_439_io_b = FullAdder_418_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_439_io_ci = FullAdder_419_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_440_io_a = FullAdder_402_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_440_io_b = FullAdder_419_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_440_io_ci = FullAdder_420_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_441_io_a = FullAdder_403_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_441_io_b = FullAdder_420_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_441_io_ci = FullAdder_421_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_442_io_a = FullAdder_404_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_442_io_b = FullAdder_421_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_442_io_ci = FullAdder_422_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_443_io_a = HalfAdder_9_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_443_io_b = FullAdder_422_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_443_io_ci = FullAdder_423_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_444_io_a = HalfAdder_10_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_444_io_b = FullAdder_423_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_444_io_ci = FullAdder_424_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_445_io_a = HalfAdder_11_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_445_io_b = FullAdder_424_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_445_io_ci = FullAdder_425_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_446_io_a = FullAdder_396_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_446_io_b = FullAdder_405_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_446_io_ci = FullAdder_426_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_447_io_a = FullAdder_381_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_447_io_b = FullAdder_397_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_447_io_ci = FullAdder_427_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_448_io_a = FullAdder_74_io_s; // @[wallaced.scala 88:18]
  assign FullAdder_448_io_b = FullAdder_278_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_448_io_ci = FullAdder_428_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_449_io_a = FullAdder_405_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_449_io_b = FullAdder_425_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_449_io_ci = FullAdder_446_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_450_io_a = FullAdder_397_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_450_io_b = FullAdder_406_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_450_io_ci = FullAdder_447_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_451_io_a = FullAdder_278_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_451_io_b = FullAdder_328_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_451_io_ci = FullAdder_448_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_452_io_a = FullAdder_328_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_452_io_b = FullAdder_360_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_452_io_ci = FullAdder_451_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_453_io_a = FullAdder_406_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_453_io_b = FullAdder_426_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_453_io_ci = FullAdder_450_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_454_io_a = FullAdder_360_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_454_io_b = FullAdder_382_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_454_io_ci = FullAdder_452_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_455_io_a = FullAdder_382_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_455_io_b = FullAdder_398_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_455_io_ci = FullAdder_454_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_456_io_a = FullAdder_398_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_456_io_b = FullAdder_407_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_456_io_ci = FullAdder_455_io_co; // @[wallaced.scala 90:19]
  assign FullAdder_457_io_a = FullAdder_407_io_co; // @[wallaced.scala 88:18]
  assign FullAdder_457_io_b = FullAdder_427_io_s; // @[wallaced.scala 89:18]
  assign FullAdder_457_io_ci = FullAdder_456_io_co; // @[wallaced.scala 90:19]
endmodule
module Black(
  input   io_i_pj,
  input   io_i_gj,
  input   io_i_pk,
  input   io_i_gk,
  output  io_o_g,
  output  io_o_p
);
  wire  _T = io_i_gj & io_i_pk; // @[pg.scala 26:32]
  assign io_o_g = io_i_gk | _T; // @[pg.scala 26:10]
  assign io_o_p = io_i_pk & io_i_pj; // @[pg.scala 27:10]
endmodule
module PPAdder(
  input         clock,
  input         reset,
  input  [31:0] io_augend,
  input  [31:0] io_addend,
  output [31:0] io_outs
);
  wire  PG_io_a; // @[ppadder.scala 35:20]
  wire  PG_io_b; // @[ppadder.scala 35:20]
  wire  PG_io_s; // @[ppadder.scala 35:20]
  wire  PG_io_co; // @[ppadder.scala 35:20]
  wire  PG_1_io_a; // @[ppadder.scala 35:20]
  wire  PG_1_io_b; // @[ppadder.scala 35:20]
  wire  PG_1_io_s; // @[ppadder.scala 35:20]
  wire  PG_1_io_co; // @[ppadder.scala 35:20]
  wire  PG_2_io_a; // @[ppadder.scala 35:20]
  wire  PG_2_io_b; // @[ppadder.scala 35:20]
  wire  PG_2_io_s; // @[ppadder.scala 35:20]
  wire  PG_2_io_co; // @[ppadder.scala 35:20]
  wire  PG_3_io_a; // @[ppadder.scala 35:20]
  wire  PG_3_io_b; // @[ppadder.scala 35:20]
  wire  PG_3_io_s; // @[ppadder.scala 35:20]
  wire  PG_3_io_co; // @[ppadder.scala 35:20]
  wire  PG_4_io_a; // @[ppadder.scala 35:20]
  wire  PG_4_io_b; // @[ppadder.scala 35:20]
  wire  PG_4_io_s; // @[ppadder.scala 35:20]
  wire  PG_4_io_co; // @[ppadder.scala 35:20]
  wire  PG_5_io_a; // @[ppadder.scala 35:20]
  wire  PG_5_io_b; // @[ppadder.scala 35:20]
  wire  PG_5_io_s; // @[ppadder.scala 35:20]
  wire  PG_5_io_co; // @[ppadder.scala 35:20]
  wire  PG_6_io_a; // @[ppadder.scala 35:20]
  wire  PG_6_io_b; // @[ppadder.scala 35:20]
  wire  PG_6_io_s; // @[ppadder.scala 35:20]
  wire  PG_6_io_co; // @[ppadder.scala 35:20]
  wire  PG_7_io_a; // @[ppadder.scala 35:20]
  wire  PG_7_io_b; // @[ppadder.scala 35:20]
  wire  PG_7_io_s; // @[ppadder.scala 35:20]
  wire  PG_7_io_co; // @[ppadder.scala 35:20]
  wire  PG_8_io_a; // @[ppadder.scala 35:20]
  wire  PG_8_io_b; // @[ppadder.scala 35:20]
  wire  PG_8_io_s; // @[ppadder.scala 35:20]
  wire  PG_8_io_co; // @[ppadder.scala 35:20]
  wire  PG_9_io_a; // @[ppadder.scala 35:20]
  wire  PG_9_io_b; // @[ppadder.scala 35:20]
  wire  PG_9_io_s; // @[ppadder.scala 35:20]
  wire  PG_9_io_co; // @[ppadder.scala 35:20]
  wire  PG_10_io_a; // @[ppadder.scala 35:20]
  wire  PG_10_io_b; // @[ppadder.scala 35:20]
  wire  PG_10_io_s; // @[ppadder.scala 35:20]
  wire  PG_10_io_co; // @[ppadder.scala 35:20]
  wire  PG_11_io_a; // @[ppadder.scala 35:20]
  wire  PG_11_io_b; // @[ppadder.scala 35:20]
  wire  PG_11_io_s; // @[ppadder.scala 35:20]
  wire  PG_11_io_co; // @[ppadder.scala 35:20]
  wire  PG_12_io_a; // @[ppadder.scala 35:20]
  wire  PG_12_io_b; // @[ppadder.scala 35:20]
  wire  PG_12_io_s; // @[ppadder.scala 35:20]
  wire  PG_12_io_co; // @[ppadder.scala 35:20]
  wire  PG_13_io_a; // @[ppadder.scala 35:20]
  wire  PG_13_io_b; // @[ppadder.scala 35:20]
  wire  PG_13_io_s; // @[ppadder.scala 35:20]
  wire  PG_13_io_co; // @[ppadder.scala 35:20]
  wire  PG_14_io_a; // @[ppadder.scala 35:20]
  wire  PG_14_io_b; // @[ppadder.scala 35:20]
  wire  PG_14_io_s; // @[ppadder.scala 35:20]
  wire  PG_14_io_co; // @[ppadder.scala 35:20]
  wire  PG_15_io_a; // @[ppadder.scala 35:20]
  wire  PG_15_io_b; // @[ppadder.scala 35:20]
  wire  PG_15_io_s; // @[ppadder.scala 35:20]
  wire  PG_15_io_co; // @[ppadder.scala 35:20]
  wire  PG_16_io_a; // @[ppadder.scala 35:20]
  wire  PG_16_io_b; // @[ppadder.scala 35:20]
  wire  PG_16_io_s; // @[ppadder.scala 35:20]
  wire  PG_16_io_co; // @[ppadder.scala 35:20]
  wire  PG_17_io_a; // @[ppadder.scala 35:20]
  wire  PG_17_io_b; // @[ppadder.scala 35:20]
  wire  PG_17_io_s; // @[ppadder.scala 35:20]
  wire  PG_17_io_co; // @[ppadder.scala 35:20]
  wire  PG_18_io_a; // @[ppadder.scala 35:20]
  wire  PG_18_io_b; // @[ppadder.scala 35:20]
  wire  PG_18_io_s; // @[ppadder.scala 35:20]
  wire  PG_18_io_co; // @[ppadder.scala 35:20]
  wire  PG_19_io_a; // @[ppadder.scala 35:20]
  wire  PG_19_io_b; // @[ppadder.scala 35:20]
  wire  PG_19_io_s; // @[ppadder.scala 35:20]
  wire  PG_19_io_co; // @[ppadder.scala 35:20]
  wire  PG_20_io_a; // @[ppadder.scala 35:20]
  wire  PG_20_io_b; // @[ppadder.scala 35:20]
  wire  PG_20_io_s; // @[ppadder.scala 35:20]
  wire  PG_20_io_co; // @[ppadder.scala 35:20]
  wire  PG_21_io_a; // @[ppadder.scala 35:20]
  wire  PG_21_io_b; // @[ppadder.scala 35:20]
  wire  PG_21_io_s; // @[ppadder.scala 35:20]
  wire  PG_21_io_co; // @[ppadder.scala 35:20]
  wire  PG_22_io_a; // @[ppadder.scala 35:20]
  wire  PG_22_io_b; // @[ppadder.scala 35:20]
  wire  PG_22_io_s; // @[ppadder.scala 35:20]
  wire  PG_22_io_co; // @[ppadder.scala 35:20]
  wire  PG_23_io_a; // @[ppadder.scala 35:20]
  wire  PG_23_io_b; // @[ppadder.scala 35:20]
  wire  PG_23_io_s; // @[ppadder.scala 35:20]
  wire  PG_23_io_co; // @[ppadder.scala 35:20]
  wire  PG_24_io_a; // @[ppadder.scala 35:20]
  wire  PG_24_io_b; // @[ppadder.scala 35:20]
  wire  PG_24_io_s; // @[ppadder.scala 35:20]
  wire  PG_24_io_co; // @[ppadder.scala 35:20]
  wire  PG_25_io_a; // @[ppadder.scala 35:20]
  wire  PG_25_io_b; // @[ppadder.scala 35:20]
  wire  PG_25_io_s; // @[ppadder.scala 35:20]
  wire  PG_25_io_co; // @[ppadder.scala 35:20]
  wire  PG_26_io_a; // @[ppadder.scala 35:20]
  wire  PG_26_io_b; // @[ppadder.scala 35:20]
  wire  PG_26_io_s; // @[ppadder.scala 35:20]
  wire  PG_26_io_co; // @[ppadder.scala 35:20]
  wire  PG_27_io_a; // @[ppadder.scala 35:20]
  wire  PG_27_io_b; // @[ppadder.scala 35:20]
  wire  PG_27_io_s; // @[ppadder.scala 35:20]
  wire  PG_27_io_co; // @[ppadder.scala 35:20]
  wire  PG_28_io_a; // @[ppadder.scala 35:20]
  wire  PG_28_io_b; // @[ppadder.scala 35:20]
  wire  PG_28_io_s; // @[ppadder.scala 35:20]
  wire  PG_28_io_co; // @[ppadder.scala 35:20]
  wire  PG_29_io_a; // @[ppadder.scala 35:20]
  wire  PG_29_io_b; // @[ppadder.scala 35:20]
  wire  PG_29_io_s; // @[ppadder.scala 35:20]
  wire  PG_29_io_co; // @[ppadder.scala 35:20]
  wire  PG_30_io_a; // @[ppadder.scala 35:20]
  wire  PG_30_io_b; // @[ppadder.scala 35:20]
  wire  PG_30_io_s; // @[ppadder.scala 35:20]
  wire  PG_30_io_co; // @[ppadder.scala 35:20]
  wire  PG_31_io_a; // @[ppadder.scala 35:20]
  wire  PG_31_io_b; // @[ppadder.scala 35:20]
  wire  PG_31_io_s; // @[ppadder.scala 35:20]
  wire  PG_31_io_co; // @[ppadder.scala 35:20]
  wire  Black_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_1_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_1_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_2_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_2_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_3_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_3_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_4_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_4_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_5_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_5_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_6_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_6_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_7_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_7_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_8_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_8_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_9_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_9_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_10_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_10_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_11_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_11_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_12_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_12_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_13_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_13_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_14_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_14_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_15_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_15_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_16_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_16_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_17_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_17_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_18_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_18_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_19_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_19_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_20_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_20_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_21_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_21_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_22_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_22_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_23_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_23_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_24_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_24_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_25_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_25_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_26_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_26_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_27_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_27_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_28_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_28_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_29_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_29_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_30_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_30_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_31_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_31_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_32_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_32_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_33_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_33_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_34_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_34_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_35_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_35_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_36_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_36_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_37_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_37_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_38_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_38_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_39_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_39_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_40_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_40_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_41_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_41_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_42_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_42_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_43_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_43_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_44_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_44_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_45_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_45_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_46_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_46_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_47_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_47_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_48_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_48_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_49_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_49_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_50_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_50_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_51_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_51_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_52_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_52_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_53_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_53_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_54_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_54_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_55_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_55_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_56_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_56_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_57_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_57_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_58_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_58_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_59_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_59_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_60_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_60_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_61_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_61_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_62_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_62_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_62_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_62_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_62_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_62_io_o_p; // @[ppadder.scala 62:23]
  wire  res_0 = PG_io_s; // @[ppadder.scala 76:40]
  wire  _T_66 = ~reset; // @[ppadder.scala 77:9]
  wire  res_1 = PG_1_io_s ^ PG_io_co; // @[ppadder.scala 80:43]
  wire  res_2 = PG_2_io_s ^ Black_32_io_o_g; // @[ppadder.scala 80:43]
  wire  res_3 = PG_3_io_s ^ Black_61_io_o_g; // @[ppadder.scala 80:43]
  wire  res_4 = PG_4_io_s ^ Black_33_io_o_g; // @[ppadder.scala 80:43]
  wire  res_5 = PG_5_io_s ^ Black_59_io_o_g; // @[ppadder.scala 80:43]
  wire  res_6 = PG_6_io_s ^ Black_60_io_o_g; // @[ppadder.scala 80:43]
  wire  res_7 = PG_7_io_s ^ Black_34_io_o_g; // @[ppadder.scala 80:43]
  wire  res_8 = PG_8_io_s ^ Black_58_io_o_g; // @[ppadder.scala 80:43]
  wire  res_9 = PG_9_io_s ^ Black_57_io_o_g; // @[ppadder.scala 80:43]
  wire  res_10 = PG_10_io_s ^ Black_55_io_o_g; // @[ppadder.scala 80:43]
  wire  res_11 = PG_11_io_s ^ Black_56_io_o_g; // @[ppadder.scala 80:43]
  wire  res_12 = PG_12_io_s ^ Black_35_io_o_g; // @[ppadder.scala 80:43]
  wire  res_13 = PG_13_io_s ^ Black_54_io_o_g; // @[ppadder.scala 80:43]
  wire  res_14 = PG_14_io_s ^ Black_53_io_o_g; // @[ppadder.scala 80:43]
  wire  res_15 = PG_15_io_s ^ Black_52_io_o_g; // @[ppadder.scala 80:43]
  wire  res_16 = PG_16_io_s ^ Black_51_io_o_g; // @[ppadder.scala 80:43]
  wire  res_17 = PG_17_io_s ^ Black_36_io_o_g; // @[ppadder.scala 80:43]
  wire  res_18 = PG_18_io_s ^ Black_50_io_o_g; // @[ppadder.scala 80:43]
  wire  res_19 = PG_19_io_s ^ Black_49_io_o_g; // @[ppadder.scala 80:43]
  wire  res_20 = PG_20_io_s ^ Black_48_io_o_g; // @[ppadder.scala 80:43]
  wire  res_21 = PG_21_io_s ^ Black_47_io_o_g; // @[ppadder.scala 80:43]
  wire  res_22 = PG_22_io_s ^ Black_46_io_o_g; // @[ppadder.scala 80:43]
  wire  res_23 = PG_23_io_s ^ Black_45_io_o_g; // @[ppadder.scala 80:43]
  wire  res_24 = PG_24_io_s ^ Black_44_io_o_g; // @[ppadder.scala 80:43]
  wire  res_25 = PG_25_io_s ^ Black_43_io_o_g; // @[ppadder.scala 80:43]
  wire  res_26 = PG_26_io_s ^ Black_42_io_o_g; // @[ppadder.scala 80:43]
  wire  res_27 = PG_27_io_s ^ Black_41_io_o_g; // @[ppadder.scala 80:43]
  wire  res_28 = PG_28_io_s ^ Black_40_io_o_g; // @[ppadder.scala 80:43]
  wire  res_29 = PG_29_io_s ^ Black_39_io_o_g; // @[ppadder.scala 80:43]
  wire  res_30 = PG_30_io_s ^ Black_38_io_o_g; // @[ppadder.scala 80:43]
  wire  res_31 = PG_31_io_s ^ Black_37_io_o_g; // @[ppadder.scala 80:43]
  wire [9:0] _T_106 = {res_31,res_30,res_29,res_28,res_27,res_26,res_25,res_24,res_23,res_22}; // @[Cat.scala 29:58]
  wire [18:0] _T_115 = {_T_106,res_21,res_20,res_19,res_18,res_17,res_16,res_15,res_14,res_13}; // @[Cat.scala 29:58]
  wire [27:0] _T_124 = {_T_115,res_12,res_11,res_10,res_9,res_8,res_7,res_6,res_5,res_4}; // @[Cat.scala 29:58]
  wire [30:0] _T_127 = {_T_124,res_3,res_2,res_1}; // @[Cat.scala 29:58]
  HalfAdder PG ( // @[ppadder.scala 35:20]
    .io_a(PG_io_a),
    .io_b(PG_io_b),
    .io_s(PG_io_s),
    .io_co(PG_io_co)
  );
  HalfAdder PG_1 ( // @[ppadder.scala 35:20]
    .io_a(PG_1_io_a),
    .io_b(PG_1_io_b),
    .io_s(PG_1_io_s),
    .io_co(PG_1_io_co)
  );
  HalfAdder PG_2 ( // @[ppadder.scala 35:20]
    .io_a(PG_2_io_a),
    .io_b(PG_2_io_b),
    .io_s(PG_2_io_s),
    .io_co(PG_2_io_co)
  );
  HalfAdder PG_3 ( // @[ppadder.scala 35:20]
    .io_a(PG_3_io_a),
    .io_b(PG_3_io_b),
    .io_s(PG_3_io_s),
    .io_co(PG_3_io_co)
  );
  HalfAdder PG_4 ( // @[ppadder.scala 35:20]
    .io_a(PG_4_io_a),
    .io_b(PG_4_io_b),
    .io_s(PG_4_io_s),
    .io_co(PG_4_io_co)
  );
  HalfAdder PG_5 ( // @[ppadder.scala 35:20]
    .io_a(PG_5_io_a),
    .io_b(PG_5_io_b),
    .io_s(PG_5_io_s),
    .io_co(PG_5_io_co)
  );
  HalfAdder PG_6 ( // @[ppadder.scala 35:20]
    .io_a(PG_6_io_a),
    .io_b(PG_6_io_b),
    .io_s(PG_6_io_s),
    .io_co(PG_6_io_co)
  );
  HalfAdder PG_7 ( // @[ppadder.scala 35:20]
    .io_a(PG_7_io_a),
    .io_b(PG_7_io_b),
    .io_s(PG_7_io_s),
    .io_co(PG_7_io_co)
  );
  HalfAdder PG_8 ( // @[ppadder.scala 35:20]
    .io_a(PG_8_io_a),
    .io_b(PG_8_io_b),
    .io_s(PG_8_io_s),
    .io_co(PG_8_io_co)
  );
  HalfAdder PG_9 ( // @[ppadder.scala 35:20]
    .io_a(PG_9_io_a),
    .io_b(PG_9_io_b),
    .io_s(PG_9_io_s),
    .io_co(PG_9_io_co)
  );
  HalfAdder PG_10 ( // @[ppadder.scala 35:20]
    .io_a(PG_10_io_a),
    .io_b(PG_10_io_b),
    .io_s(PG_10_io_s),
    .io_co(PG_10_io_co)
  );
  HalfAdder PG_11 ( // @[ppadder.scala 35:20]
    .io_a(PG_11_io_a),
    .io_b(PG_11_io_b),
    .io_s(PG_11_io_s),
    .io_co(PG_11_io_co)
  );
  HalfAdder PG_12 ( // @[ppadder.scala 35:20]
    .io_a(PG_12_io_a),
    .io_b(PG_12_io_b),
    .io_s(PG_12_io_s),
    .io_co(PG_12_io_co)
  );
  HalfAdder PG_13 ( // @[ppadder.scala 35:20]
    .io_a(PG_13_io_a),
    .io_b(PG_13_io_b),
    .io_s(PG_13_io_s),
    .io_co(PG_13_io_co)
  );
  HalfAdder PG_14 ( // @[ppadder.scala 35:20]
    .io_a(PG_14_io_a),
    .io_b(PG_14_io_b),
    .io_s(PG_14_io_s),
    .io_co(PG_14_io_co)
  );
  HalfAdder PG_15 ( // @[ppadder.scala 35:20]
    .io_a(PG_15_io_a),
    .io_b(PG_15_io_b),
    .io_s(PG_15_io_s),
    .io_co(PG_15_io_co)
  );
  HalfAdder PG_16 ( // @[ppadder.scala 35:20]
    .io_a(PG_16_io_a),
    .io_b(PG_16_io_b),
    .io_s(PG_16_io_s),
    .io_co(PG_16_io_co)
  );
  HalfAdder PG_17 ( // @[ppadder.scala 35:20]
    .io_a(PG_17_io_a),
    .io_b(PG_17_io_b),
    .io_s(PG_17_io_s),
    .io_co(PG_17_io_co)
  );
  HalfAdder PG_18 ( // @[ppadder.scala 35:20]
    .io_a(PG_18_io_a),
    .io_b(PG_18_io_b),
    .io_s(PG_18_io_s),
    .io_co(PG_18_io_co)
  );
  HalfAdder PG_19 ( // @[ppadder.scala 35:20]
    .io_a(PG_19_io_a),
    .io_b(PG_19_io_b),
    .io_s(PG_19_io_s),
    .io_co(PG_19_io_co)
  );
  HalfAdder PG_20 ( // @[ppadder.scala 35:20]
    .io_a(PG_20_io_a),
    .io_b(PG_20_io_b),
    .io_s(PG_20_io_s),
    .io_co(PG_20_io_co)
  );
  HalfAdder PG_21 ( // @[ppadder.scala 35:20]
    .io_a(PG_21_io_a),
    .io_b(PG_21_io_b),
    .io_s(PG_21_io_s),
    .io_co(PG_21_io_co)
  );
  HalfAdder PG_22 ( // @[ppadder.scala 35:20]
    .io_a(PG_22_io_a),
    .io_b(PG_22_io_b),
    .io_s(PG_22_io_s),
    .io_co(PG_22_io_co)
  );
  HalfAdder PG_23 ( // @[ppadder.scala 35:20]
    .io_a(PG_23_io_a),
    .io_b(PG_23_io_b),
    .io_s(PG_23_io_s),
    .io_co(PG_23_io_co)
  );
  HalfAdder PG_24 ( // @[ppadder.scala 35:20]
    .io_a(PG_24_io_a),
    .io_b(PG_24_io_b),
    .io_s(PG_24_io_s),
    .io_co(PG_24_io_co)
  );
  HalfAdder PG_25 ( // @[ppadder.scala 35:20]
    .io_a(PG_25_io_a),
    .io_b(PG_25_io_b),
    .io_s(PG_25_io_s),
    .io_co(PG_25_io_co)
  );
  HalfAdder PG_26 ( // @[ppadder.scala 35:20]
    .io_a(PG_26_io_a),
    .io_b(PG_26_io_b),
    .io_s(PG_26_io_s),
    .io_co(PG_26_io_co)
  );
  HalfAdder PG_27 ( // @[ppadder.scala 35:20]
    .io_a(PG_27_io_a),
    .io_b(PG_27_io_b),
    .io_s(PG_27_io_s),
    .io_co(PG_27_io_co)
  );
  HalfAdder PG_28 ( // @[ppadder.scala 35:20]
    .io_a(PG_28_io_a),
    .io_b(PG_28_io_b),
    .io_s(PG_28_io_s),
    .io_co(PG_28_io_co)
  );
  HalfAdder PG_29 ( // @[ppadder.scala 35:20]
    .io_a(PG_29_io_a),
    .io_b(PG_29_io_b),
    .io_s(PG_29_io_s),
    .io_co(PG_29_io_co)
  );
  HalfAdder PG_30 ( // @[ppadder.scala 35:20]
    .io_a(PG_30_io_a),
    .io_b(PG_30_io_b),
    .io_s(PG_30_io_s),
    .io_co(PG_30_io_co)
  );
  HalfAdder PG_31 ( // @[ppadder.scala 35:20]
    .io_a(PG_31_io_a),
    .io_b(PG_31_io_b),
    .io_s(PG_31_io_s),
    .io_co(PG_31_io_co)
  );
  Black Black ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_io_i_pj),
    .io_i_gj(Black_io_i_gj),
    .io_i_pk(Black_io_i_pk),
    .io_i_gk(Black_io_i_gk),
    .io_o_g(Black_io_o_g),
    .io_o_p(Black_io_o_p)
  );
  Black Black_1 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_1_io_i_pj),
    .io_i_gj(Black_1_io_i_gj),
    .io_i_pk(Black_1_io_i_pk),
    .io_i_gk(Black_1_io_i_gk),
    .io_o_g(Black_1_io_o_g),
    .io_o_p(Black_1_io_o_p)
  );
  Black Black_2 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_2_io_i_pj),
    .io_i_gj(Black_2_io_i_gj),
    .io_i_pk(Black_2_io_i_pk),
    .io_i_gk(Black_2_io_i_gk),
    .io_o_g(Black_2_io_o_g),
    .io_o_p(Black_2_io_o_p)
  );
  Black Black_3 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_3_io_i_pj),
    .io_i_gj(Black_3_io_i_gj),
    .io_i_pk(Black_3_io_i_pk),
    .io_i_gk(Black_3_io_i_gk),
    .io_o_g(Black_3_io_o_g),
    .io_o_p(Black_3_io_o_p)
  );
  Black Black_4 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_4_io_i_pj),
    .io_i_gj(Black_4_io_i_gj),
    .io_i_pk(Black_4_io_i_pk),
    .io_i_gk(Black_4_io_i_gk),
    .io_o_g(Black_4_io_o_g),
    .io_o_p(Black_4_io_o_p)
  );
  Black Black_5 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_5_io_i_pj),
    .io_i_gj(Black_5_io_i_gj),
    .io_i_pk(Black_5_io_i_pk),
    .io_i_gk(Black_5_io_i_gk),
    .io_o_g(Black_5_io_o_g),
    .io_o_p(Black_5_io_o_p)
  );
  Black Black_6 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_6_io_i_pj),
    .io_i_gj(Black_6_io_i_gj),
    .io_i_pk(Black_6_io_i_pk),
    .io_i_gk(Black_6_io_i_gk),
    .io_o_g(Black_6_io_o_g),
    .io_o_p(Black_6_io_o_p)
  );
  Black Black_7 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_7_io_i_pj),
    .io_i_gj(Black_7_io_i_gj),
    .io_i_pk(Black_7_io_i_pk),
    .io_i_gk(Black_7_io_i_gk),
    .io_o_g(Black_7_io_o_g),
    .io_o_p(Black_7_io_o_p)
  );
  Black Black_8 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_8_io_i_pj),
    .io_i_gj(Black_8_io_i_gj),
    .io_i_pk(Black_8_io_i_pk),
    .io_i_gk(Black_8_io_i_gk),
    .io_o_g(Black_8_io_o_g),
    .io_o_p(Black_8_io_o_p)
  );
  Black Black_9 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_9_io_i_pj),
    .io_i_gj(Black_9_io_i_gj),
    .io_i_pk(Black_9_io_i_pk),
    .io_i_gk(Black_9_io_i_gk),
    .io_o_g(Black_9_io_o_g),
    .io_o_p(Black_9_io_o_p)
  );
  Black Black_10 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_10_io_i_pj),
    .io_i_gj(Black_10_io_i_gj),
    .io_i_pk(Black_10_io_i_pk),
    .io_i_gk(Black_10_io_i_gk),
    .io_o_g(Black_10_io_o_g),
    .io_o_p(Black_10_io_o_p)
  );
  Black Black_11 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_11_io_i_pj),
    .io_i_gj(Black_11_io_i_gj),
    .io_i_pk(Black_11_io_i_pk),
    .io_i_gk(Black_11_io_i_gk),
    .io_o_g(Black_11_io_o_g),
    .io_o_p(Black_11_io_o_p)
  );
  Black Black_12 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_12_io_i_pj),
    .io_i_gj(Black_12_io_i_gj),
    .io_i_pk(Black_12_io_i_pk),
    .io_i_gk(Black_12_io_i_gk),
    .io_o_g(Black_12_io_o_g),
    .io_o_p(Black_12_io_o_p)
  );
  Black Black_13 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_13_io_i_pj),
    .io_i_gj(Black_13_io_i_gj),
    .io_i_pk(Black_13_io_i_pk),
    .io_i_gk(Black_13_io_i_gk),
    .io_o_g(Black_13_io_o_g),
    .io_o_p(Black_13_io_o_p)
  );
  Black Black_14 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_14_io_i_pj),
    .io_i_gj(Black_14_io_i_gj),
    .io_i_pk(Black_14_io_i_pk),
    .io_i_gk(Black_14_io_i_gk),
    .io_o_g(Black_14_io_o_g),
    .io_o_p(Black_14_io_o_p)
  );
  Black Black_15 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_15_io_i_pj),
    .io_i_gj(Black_15_io_i_gj),
    .io_i_pk(Black_15_io_i_pk),
    .io_i_gk(Black_15_io_i_gk),
    .io_o_g(Black_15_io_o_g),
    .io_o_p(Black_15_io_o_p)
  );
  Black Black_16 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_16_io_i_pj),
    .io_i_gj(Black_16_io_i_gj),
    .io_i_pk(Black_16_io_i_pk),
    .io_i_gk(Black_16_io_i_gk),
    .io_o_g(Black_16_io_o_g),
    .io_o_p(Black_16_io_o_p)
  );
  Black Black_17 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_17_io_i_pj),
    .io_i_gj(Black_17_io_i_gj),
    .io_i_pk(Black_17_io_i_pk),
    .io_i_gk(Black_17_io_i_gk),
    .io_o_g(Black_17_io_o_g),
    .io_o_p(Black_17_io_o_p)
  );
  Black Black_18 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_18_io_i_pj),
    .io_i_gj(Black_18_io_i_gj),
    .io_i_pk(Black_18_io_i_pk),
    .io_i_gk(Black_18_io_i_gk),
    .io_o_g(Black_18_io_o_g),
    .io_o_p(Black_18_io_o_p)
  );
  Black Black_19 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_19_io_i_pj),
    .io_i_gj(Black_19_io_i_gj),
    .io_i_pk(Black_19_io_i_pk),
    .io_i_gk(Black_19_io_i_gk),
    .io_o_g(Black_19_io_o_g),
    .io_o_p(Black_19_io_o_p)
  );
  Black Black_20 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_20_io_i_pj),
    .io_i_gj(Black_20_io_i_gj),
    .io_i_pk(Black_20_io_i_pk),
    .io_i_gk(Black_20_io_i_gk),
    .io_o_g(Black_20_io_o_g),
    .io_o_p(Black_20_io_o_p)
  );
  Black Black_21 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_21_io_i_pj),
    .io_i_gj(Black_21_io_i_gj),
    .io_i_pk(Black_21_io_i_pk),
    .io_i_gk(Black_21_io_i_gk),
    .io_o_g(Black_21_io_o_g),
    .io_o_p(Black_21_io_o_p)
  );
  Black Black_22 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_22_io_i_pj),
    .io_i_gj(Black_22_io_i_gj),
    .io_i_pk(Black_22_io_i_pk),
    .io_i_gk(Black_22_io_i_gk),
    .io_o_g(Black_22_io_o_g),
    .io_o_p(Black_22_io_o_p)
  );
  Black Black_23 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_23_io_i_pj),
    .io_i_gj(Black_23_io_i_gj),
    .io_i_pk(Black_23_io_i_pk),
    .io_i_gk(Black_23_io_i_gk),
    .io_o_g(Black_23_io_o_g),
    .io_o_p(Black_23_io_o_p)
  );
  Black Black_24 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_24_io_i_pj),
    .io_i_gj(Black_24_io_i_gj),
    .io_i_pk(Black_24_io_i_pk),
    .io_i_gk(Black_24_io_i_gk),
    .io_o_g(Black_24_io_o_g),
    .io_o_p(Black_24_io_o_p)
  );
  Black Black_25 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_25_io_i_pj),
    .io_i_gj(Black_25_io_i_gj),
    .io_i_pk(Black_25_io_i_pk),
    .io_i_gk(Black_25_io_i_gk),
    .io_o_g(Black_25_io_o_g),
    .io_o_p(Black_25_io_o_p)
  );
  Black Black_26 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_26_io_i_pj),
    .io_i_gj(Black_26_io_i_gj),
    .io_i_pk(Black_26_io_i_pk),
    .io_i_gk(Black_26_io_i_gk),
    .io_o_g(Black_26_io_o_g),
    .io_o_p(Black_26_io_o_p)
  );
  Black Black_27 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_27_io_i_pj),
    .io_i_gj(Black_27_io_i_gj),
    .io_i_pk(Black_27_io_i_pk),
    .io_i_gk(Black_27_io_i_gk),
    .io_o_g(Black_27_io_o_g),
    .io_o_p(Black_27_io_o_p)
  );
  Black Black_28 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_28_io_i_pj),
    .io_i_gj(Black_28_io_i_gj),
    .io_i_pk(Black_28_io_i_pk),
    .io_i_gk(Black_28_io_i_gk),
    .io_o_g(Black_28_io_o_g),
    .io_o_p(Black_28_io_o_p)
  );
  Black Black_29 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_29_io_i_pj),
    .io_i_gj(Black_29_io_i_gj),
    .io_i_pk(Black_29_io_i_pk),
    .io_i_gk(Black_29_io_i_gk),
    .io_o_g(Black_29_io_o_g),
    .io_o_p(Black_29_io_o_p)
  );
  Black Black_30 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_30_io_i_pj),
    .io_i_gj(Black_30_io_i_gj),
    .io_i_pk(Black_30_io_i_pk),
    .io_i_gk(Black_30_io_i_gk),
    .io_o_g(Black_30_io_o_g),
    .io_o_p(Black_30_io_o_p)
  );
  Black Black_31 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_31_io_i_pj),
    .io_i_gj(Black_31_io_i_gj),
    .io_i_pk(Black_31_io_i_pk),
    .io_i_gk(Black_31_io_i_gk),
    .io_o_g(Black_31_io_o_g),
    .io_o_p(Black_31_io_o_p)
  );
  Black Black_32 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_32_io_i_pj),
    .io_i_gj(Black_32_io_i_gj),
    .io_i_pk(Black_32_io_i_pk),
    .io_i_gk(Black_32_io_i_gk),
    .io_o_g(Black_32_io_o_g),
    .io_o_p(Black_32_io_o_p)
  );
  Black Black_33 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_33_io_i_pj),
    .io_i_gj(Black_33_io_i_gj),
    .io_i_pk(Black_33_io_i_pk),
    .io_i_gk(Black_33_io_i_gk),
    .io_o_g(Black_33_io_o_g),
    .io_o_p(Black_33_io_o_p)
  );
  Black Black_34 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_34_io_i_pj),
    .io_i_gj(Black_34_io_i_gj),
    .io_i_pk(Black_34_io_i_pk),
    .io_i_gk(Black_34_io_i_gk),
    .io_o_g(Black_34_io_o_g),
    .io_o_p(Black_34_io_o_p)
  );
  Black Black_35 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_35_io_i_pj),
    .io_i_gj(Black_35_io_i_gj),
    .io_i_pk(Black_35_io_i_pk),
    .io_i_gk(Black_35_io_i_gk),
    .io_o_g(Black_35_io_o_g),
    .io_o_p(Black_35_io_o_p)
  );
  Black Black_36 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_36_io_i_pj),
    .io_i_gj(Black_36_io_i_gj),
    .io_i_pk(Black_36_io_i_pk),
    .io_i_gk(Black_36_io_i_gk),
    .io_o_g(Black_36_io_o_g),
    .io_o_p(Black_36_io_o_p)
  );
  Black Black_37 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_37_io_i_pj),
    .io_i_gj(Black_37_io_i_gj),
    .io_i_pk(Black_37_io_i_pk),
    .io_i_gk(Black_37_io_i_gk),
    .io_o_g(Black_37_io_o_g),
    .io_o_p(Black_37_io_o_p)
  );
  Black Black_38 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_38_io_i_pj),
    .io_i_gj(Black_38_io_i_gj),
    .io_i_pk(Black_38_io_i_pk),
    .io_i_gk(Black_38_io_i_gk),
    .io_o_g(Black_38_io_o_g),
    .io_o_p(Black_38_io_o_p)
  );
  Black Black_39 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_39_io_i_pj),
    .io_i_gj(Black_39_io_i_gj),
    .io_i_pk(Black_39_io_i_pk),
    .io_i_gk(Black_39_io_i_gk),
    .io_o_g(Black_39_io_o_g),
    .io_o_p(Black_39_io_o_p)
  );
  Black Black_40 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_40_io_i_pj),
    .io_i_gj(Black_40_io_i_gj),
    .io_i_pk(Black_40_io_i_pk),
    .io_i_gk(Black_40_io_i_gk),
    .io_o_g(Black_40_io_o_g),
    .io_o_p(Black_40_io_o_p)
  );
  Black Black_41 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_41_io_i_pj),
    .io_i_gj(Black_41_io_i_gj),
    .io_i_pk(Black_41_io_i_pk),
    .io_i_gk(Black_41_io_i_gk),
    .io_o_g(Black_41_io_o_g),
    .io_o_p(Black_41_io_o_p)
  );
  Black Black_42 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_42_io_i_pj),
    .io_i_gj(Black_42_io_i_gj),
    .io_i_pk(Black_42_io_i_pk),
    .io_i_gk(Black_42_io_i_gk),
    .io_o_g(Black_42_io_o_g),
    .io_o_p(Black_42_io_o_p)
  );
  Black Black_43 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_43_io_i_pj),
    .io_i_gj(Black_43_io_i_gj),
    .io_i_pk(Black_43_io_i_pk),
    .io_i_gk(Black_43_io_i_gk),
    .io_o_g(Black_43_io_o_g),
    .io_o_p(Black_43_io_o_p)
  );
  Black Black_44 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_44_io_i_pj),
    .io_i_gj(Black_44_io_i_gj),
    .io_i_pk(Black_44_io_i_pk),
    .io_i_gk(Black_44_io_i_gk),
    .io_o_g(Black_44_io_o_g),
    .io_o_p(Black_44_io_o_p)
  );
  Black Black_45 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_45_io_i_pj),
    .io_i_gj(Black_45_io_i_gj),
    .io_i_pk(Black_45_io_i_pk),
    .io_i_gk(Black_45_io_i_gk),
    .io_o_g(Black_45_io_o_g),
    .io_o_p(Black_45_io_o_p)
  );
  Black Black_46 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_46_io_i_pj),
    .io_i_gj(Black_46_io_i_gj),
    .io_i_pk(Black_46_io_i_pk),
    .io_i_gk(Black_46_io_i_gk),
    .io_o_g(Black_46_io_o_g),
    .io_o_p(Black_46_io_o_p)
  );
  Black Black_47 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_47_io_i_pj),
    .io_i_gj(Black_47_io_i_gj),
    .io_i_pk(Black_47_io_i_pk),
    .io_i_gk(Black_47_io_i_gk),
    .io_o_g(Black_47_io_o_g),
    .io_o_p(Black_47_io_o_p)
  );
  Black Black_48 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_48_io_i_pj),
    .io_i_gj(Black_48_io_i_gj),
    .io_i_pk(Black_48_io_i_pk),
    .io_i_gk(Black_48_io_i_gk),
    .io_o_g(Black_48_io_o_g),
    .io_o_p(Black_48_io_o_p)
  );
  Black Black_49 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_49_io_i_pj),
    .io_i_gj(Black_49_io_i_gj),
    .io_i_pk(Black_49_io_i_pk),
    .io_i_gk(Black_49_io_i_gk),
    .io_o_g(Black_49_io_o_g),
    .io_o_p(Black_49_io_o_p)
  );
  Black Black_50 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_50_io_i_pj),
    .io_i_gj(Black_50_io_i_gj),
    .io_i_pk(Black_50_io_i_pk),
    .io_i_gk(Black_50_io_i_gk),
    .io_o_g(Black_50_io_o_g),
    .io_o_p(Black_50_io_o_p)
  );
  Black Black_51 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_51_io_i_pj),
    .io_i_gj(Black_51_io_i_gj),
    .io_i_pk(Black_51_io_i_pk),
    .io_i_gk(Black_51_io_i_gk),
    .io_o_g(Black_51_io_o_g),
    .io_o_p(Black_51_io_o_p)
  );
  Black Black_52 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_52_io_i_pj),
    .io_i_gj(Black_52_io_i_gj),
    .io_i_pk(Black_52_io_i_pk),
    .io_i_gk(Black_52_io_i_gk),
    .io_o_g(Black_52_io_o_g),
    .io_o_p(Black_52_io_o_p)
  );
  Black Black_53 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_53_io_i_pj),
    .io_i_gj(Black_53_io_i_gj),
    .io_i_pk(Black_53_io_i_pk),
    .io_i_gk(Black_53_io_i_gk),
    .io_o_g(Black_53_io_o_g),
    .io_o_p(Black_53_io_o_p)
  );
  Black Black_54 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_54_io_i_pj),
    .io_i_gj(Black_54_io_i_gj),
    .io_i_pk(Black_54_io_i_pk),
    .io_i_gk(Black_54_io_i_gk),
    .io_o_g(Black_54_io_o_g),
    .io_o_p(Black_54_io_o_p)
  );
  Black Black_55 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_55_io_i_pj),
    .io_i_gj(Black_55_io_i_gj),
    .io_i_pk(Black_55_io_i_pk),
    .io_i_gk(Black_55_io_i_gk),
    .io_o_g(Black_55_io_o_g),
    .io_o_p(Black_55_io_o_p)
  );
  Black Black_56 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_56_io_i_pj),
    .io_i_gj(Black_56_io_i_gj),
    .io_i_pk(Black_56_io_i_pk),
    .io_i_gk(Black_56_io_i_gk),
    .io_o_g(Black_56_io_o_g),
    .io_o_p(Black_56_io_o_p)
  );
  Black Black_57 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_57_io_i_pj),
    .io_i_gj(Black_57_io_i_gj),
    .io_i_pk(Black_57_io_i_pk),
    .io_i_gk(Black_57_io_i_gk),
    .io_o_g(Black_57_io_o_g),
    .io_o_p(Black_57_io_o_p)
  );
  Black Black_58 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_58_io_i_pj),
    .io_i_gj(Black_58_io_i_gj),
    .io_i_pk(Black_58_io_i_pk),
    .io_i_gk(Black_58_io_i_gk),
    .io_o_g(Black_58_io_o_g),
    .io_o_p(Black_58_io_o_p)
  );
  Black Black_59 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_59_io_i_pj),
    .io_i_gj(Black_59_io_i_gj),
    .io_i_pk(Black_59_io_i_pk),
    .io_i_gk(Black_59_io_i_gk),
    .io_o_g(Black_59_io_o_g),
    .io_o_p(Black_59_io_o_p)
  );
  Black Black_60 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_60_io_i_pj),
    .io_i_gj(Black_60_io_i_gj),
    .io_i_pk(Black_60_io_i_pk),
    .io_i_gk(Black_60_io_i_gk),
    .io_o_g(Black_60_io_o_g),
    .io_o_p(Black_60_io_o_p)
  );
  Black Black_61 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_61_io_i_pj),
    .io_i_gj(Black_61_io_i_gj),
    .io_i_pk(Black_61_io_i_pk),
    .io_i_gk(Black_61_io_i_gk),
    .io_o_g(Black_61_io_o_g),
    .io_o_p(Black_61_io_o_p)
  );
  Black Black_62 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_62_io_i_pj),
    .io_i_gj(Black_62_io_i_gj),
    .io_i_pk(Black_62_io_i_pk),
    .io_i_gk(Black_62_io_i_gk),
    .io_o_g(Black_62_io_o_g),
    .io_o_p(Black_62_io_o_p)
  );
  assign io_outs = {_T_127,res_0}; // @[ppadder.scala 84:11]
  assign PG_io_a = io_augend[0]; // @[ppadder.scala 36:15]
  assign PG_io_b = io_addend[0]; // @[ppadder.scala 37:15]
  assign PG_1_io_a = io_augend[1]; // @[ppadder.scala 36:15]
  assign PG_1_io_b = io_addend[1]; // @[ppadder.scala 37:15]
  assign PG_2_io_a = io_augend[2]; // @[ppadder.scala 36:15]
  assign PG_2_io_b = io_addend[2]; // @[ppadder.scala 37:15]
  assign PG_3_io_a = io_augend[3]; // @[ppadder.scala 36:15]
  assign PG_3_io_b = io_addend[3]; // @[ppadder.scala 37:15]
  assign PG_4_io_a = io_augend[4]; // @[ppadder.scala 36:15]
  assign PG_4_io_b = io_addend[4]; // @[ppadder.scala 37:15]
  assign PG_5_io_a = io_augend[5]; // @[ppadder.scala 36:15]
  assign PG_5_io_b = io_addend[5]; // @[ppadder.scala 37:15]
  assign PG_6_io_a = io_augend[6]; // @[ppadder.scala 36:15]
  assign PG_6_io_b = io_addend[6]; // @[ppadder.scala 37:15]
  assign PG_7_io_a = io_augend[7]; // @[ppadder.scala 36:15]
  assign PG_7_io_b = io_addend[7]; // @[ppadder.scala 37:15]
  assign PG_8_io_a = io_augend[8]; // @[ppadder.scala 36:15]
  assign PG_8_io_b = io_addend[8]; // @[ppadder.scala 37:15]
  assign PG_9_io_a = io_augend[9]; // @[ppadder.scala 36:15]
  assign PG_9_io_b = io_addend[9]; // @[ppadder.scala 37:15]
  assign PG_10_io_a = io_augend[10]; // @[ppadder.scala 36:15]
  assign PG_10_io_b = io_addend[10]; // @[ppadder.scala 37:15]
  assign PG_11_io_a = io_augend[11]; // @[ppadder.scala 36:15]
  assign PG_11_io_b = io_addend[11]; // @[ppadder.scala 37:15]
  assign PG_12_io_a = io_augend[12]; // @[ppadder.scala 36:15]
  assign PG_12_io_b = io_addend[12]; // @[ppadder.scala 37:15]
  assign PG_13_io_a = io_augend[13]; // @[ppadder.scala 36:15]
  assign PG_13_io_b = io_addend[13]; // @[ppadder.scala 37:15]
  assign PG_14_io_a = io_augend[14]; // @[ppadder.scala 36:15]
  assign PG_14_io_b = io_addend[14]; // @[ppadder.scala 37:15]
  assign PG_15_io_a = io_augend[15]; // @[ppadder.scala 36:15]
  assign PG_15_io_b = io_addend[15]; // @[ppadder.scala 37:15]
  assign PG_16_io_a = io_augend[16]; // @[ppadder.scala 36:15]
  assign PG_16_io_b = io_addend[16]; // @[ppadder.scala 37:15]
  assign PG_17_io_a = io_augend[17]; // @[ppadder.scala 36:15]
  assign PG_17_io_b = io_addend[17]; // @[ppadder.scala 37:15]
  assign PG_18_io_a = io_augend[18]; // @[ppadder.scala 36:15]
  assign PG_18_io_b = io_addend[18]; // @[ppadder.scala 37:15]
  assign PG_19_io_a = io_augend[19]; // @[ppadder.scala 36:15]
  assign PG_19_io_b = io_addend[19]; // @[ppadder.scala 37:15]
  assign PG_20_io_a = io_augend[20]; // @[ppadder.scala 36:15]
  assign PG_20_io_b = io_addend[20]; // @[ppadder.scala 37:15]
  assign PG_21_io_a = io_augend[21]; // @[ppadder.scala 36:15]
  assign PG_21_io_b = io_addend[21]; // @[ppadder.scala 37:15]
  assign PG_22_io_a = io_augend[22]; // @[ppadder.scala 36:15]
  assign PG_22_io_b = io_addend[22]; // @[ppadder.scala 37:15]
  assign PG_23_io_a = io_augend[23]; // @[ppadder.scala 36:15]
  assign PG_23_io_b = io_addend[23]; // @[ppadder.scala 37:15]
  assign PG_24_io_a = io_augend[24]; // @[ppadder.scala 36:15]
  assign PG_24_io_b = io_addend[24]; // @[ppadder.scala 37:15]
  assign PG_25_io_a = io_augend[25]; // @[ppadder.scala 36:15]
  assign PG_25_io_b = io_addend[25]; // @[ppadder.scala 37:15]
  assign PG_26_io_a = io_augend[26]; // @[ppadder.scala 36:15]
  assign PG_26_io_b = io_addend[26]; // @[ppadder.scala 37:15]
  assign PG_27_io_a = io_augend[27]; // @[ppadder.scala 36:15]
  assign PG_27_io_b = io_addend[27]; // @[ppadder.scala 37:15]
  assign PG_28_io_a = io_augend[28]; // @[ppadder.scala 36:15]
  assign PG_28_io_b = io_addend[28]; // @[ppadder.scala 37:15]
  assign PG_29_io_a = io_augend[29]; // @[ppadder.scala 36:15]
  assign PG_29_io_b = io_addend[29]; // @[ppadder.scala 37:15]
  assign PG_30_io_a = io_augend[30]; // @[ppadder.scala 36:15]
  assign PG_30_io_b = io_addend[30]; // @[ppadder.scala 37:15]
  assign PG_31_io_a = io_augend[31]; // @[ppadder.scala 36:15]
  assign PG_31_io_b = io_addend[31]; // @[ppadder.scala 37:15]
  assign Black_io_i_pj = PG_26_io_s; // @[ppadder.scala 66:19]
  assign Black_io_i_gj = PG_26_io_co; // @[ppadder.scala 65:19]
  assign Black_io_i_pk = PG_27_io_s; // @[ppadder.scala 64:19]
  assign Black_io_i_gk = PG_27_io_co; // @[ppadder.scala 63:19]
  assign Black_1_io_i_pj = Black_io_o_p; // @[ppadder.scala 66:19]
  assign Black_1_io_i_gj = Black_io_o_g; // @[ppadder.scala 65:19]
  assign Black_1_io_i_pk = PG_28_io_s; // @[ppadder.scala 64:19]
  assign Black_1_io_i_gk = PG_28_io_co; // @[ppadder.scala 63:19]
  assign Black_2_io_i_pj = Black_1_io_o_p; // @[ppadder.scala 66:19]
  assign Black_2_io_i_gj = Black_1_io_o_g; // @[ppadder.scala 65:19]
  assign Black_2_io_i_pk = PG_29_io_s; // @[ppadder.scala 64:19]
  assign Black_2_io_i_gk = PG_29_io_co; // @[ppadder.scala 63:19]
  assign Black_3_io_i_pj = Black_2_io_o_p; // @[ppadder.scala 66:19]
  assign Black_3_io_i_gj = Black_2_io_o_g; // @[ppadder.scala 65:19]
  assign Black_3_io_i_pk = PG_30_io_s; // @[ppadder.scala 64:19]
  assign Black_3_io_i_gk = PG_30_io_co; // @[ppadder.scala 63:19]
  assign Black_4_io_i_pj = PG_22_io_s; // @[ppadder.scala 66:19]
  assign Black_4_io_i_gj = PG_22_io_co; // @[ppadder.scala 65:19]
  assign Black_4_io_i_pk = PG_23_io_s; // @[ppadder.scala 64:19]
  assign Black_4_io_i_gk = PG_23_io_co; // @[ppadder.scala 63:19]
  assign Black_5_io_i_pj = Black_4_io_o_p; // @[ppadder.scala 66:19]
  assign Black_5_io_i_gj = Black_4_io_o_g; // @[ppadder.scala 65:19]
  assign Black_5_io_i_pk = PG_24_io_s; // @[ppadder.scala 64:19]
  assign Black_5_io_i_gk = PG_24_io_co; // @[ppadder.scala 63:19]
  assign Black_6_io_i_pj = Black_5_io_o_p; // @[ppadder.scala 66:19]
  assign Black_6_io_i_gj = Black_5_io_o_g; // @[ppadder.scala 65:19]
  assign Black_6_io_i_pk = PG_25_io_s; // @[ppadder.scala 64:19]
  assign Black_6_io_i_gk = PG_25_io_co; // @[ppadder.scala 63:19]
  assign Black_7_io_i_pj = PG_20_io_s; // @[ppadder.scala 66:19]
  assign Black_7_io_i_gj = PG_20_io_co; // @[ppadder.scala 65:19]
  assign Black_7_io_i_pk = PG_21_io_s; // @[ppadder.scala 64:19]
  assign Black_7_io_i_gk = PG_21_io_co; // @[ppadder.scala 63:19]
  assign Black_8_io_i_pj = PG_17_io_s; // @[ppadder.scala 66:19]
  assign Black_8_io_i_gj = PG_17_io_co; // @[ppadder.scala 65:19]
  assign Black_8_io_i_pk = PG_18_io_s; // @[ppadder.scala 64:19]
  assign Black_8_io_i_gk = PG_18_io_co; // @[ppadder.scala 63:19]
  assign Black_9_io_i_pj = Black_8_io_o_p; // @[ppadder.scala 66:19]
  assign Black_9_io_i_gj = Black_8_io_o_g; // @[ppadder.scala 65:19]
  assign Black_9_io_i_pk = PG_19_io_s; // @[ppadder.scala 64:19]
  assign Black_9_io_i_gk = PG_19_io_co; // @[ppadder.scala 63:19]
  assign Black_10_io_i_pj = Black_9_io_o_p; // @[ppadder.scala 66:19]
  assign Black_10_io_i_gj = Black_9_io_o_g; // @[ppadder.scala 65:19]
  assign Black_10_io_i_pk = Black_7_io_o_p; // @[ppadder.scala 64:19]
  assign Black_10_io_i_gk = Black_7_io_o_g; // @[ppadder.scala 63:19]
  assign Black_11_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_11_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_11_io_i_pk = Black_6_io_o_p; // @[ppadder.scala 64:19]
  assign Black_11_io_i_gk = Black_6_io_o_g; // @[ppadder.scala 63:19]
  assign Black_12_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_12_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_12_io_i_pk = Black_3_io_o_p; // @[ppadder.scala 64:19]
  assign Black_12_io_i_gk = Black_3_io_o_g; // @[ppadder.scala 63:19]
  assign Black_13_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_13_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_13_io_i_pk = Black_2_io_o_p; // @[ppadder.scala 64:19]
  assign Black_13_io_i_gk = Black_2_io_o_g; // @[ppadder.scala 63:19]
  assign Black_14_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_14_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_14_io_i_pk = Black_1_io_o_p; // @[ppadder.scala 64:19]
  assign Black_14_io_i_gk = Black_1_io_o_g; // @[ppadder.scala 63:19]
  assign Black_15_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_15_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_15_io_i_pk = Black_io_o_p; // @[ppadder.scala 64:19]
  assign Black_15_io_i_gk = Black_io_o_g; // @[ppadder.scala 63:19]
  assign Black_16_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_16_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_16_io_i_pk = PG_26_io_s; // @[ppadder.scala 64:19]
  assign Black_16_io_i_gk = PG_26_io_co; // @[ppadder.scala 63:19]
  assign Black_17_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_17_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_17_io_i_pk = Black_5_io_o_p; // @[ppadder.scala 64:19]
  assign Black_17_io_i_gk = Black_5_io_o_g; // @[ppadder.scala 63:19]
  assign Black_18_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_18_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_18_io_i_pk = Black_4_io_o_p; // @[ppadder.scala 64:19]
  assign Black_18_io_i_gk = Black_4_io_o_g; // @[ppadder.scala 63:19]
  assign Black_19_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_19_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_19_io_i_pk = PG_22_io_s; // @[ppadder.scala 64:19]
  assign Black_19_io_i_gk = PG_22_io_co; // @[ppadder.scala 63:19]
  assign Black_20_io_i_pj = Black_9_io_o_p; // @[ppadder.scala 66:19]
  assign Black_20_io_i_gj = Black_9_io_o_g; // @[ppadder.scala 65:19]
  assign Black_20_io_i_pk = PG_20_io_s; // @[ppadder.scala 64:19]
  assign Black_20_io_i_gk = PG_20_io_co; // @[ppadder.scala 63:19]
  assign Black_21_io_i_pj = PG_12_io_s; // @[ppadder.scala 66:19]
  assign Black_21_io_i_gj = PG_12_io_co; // @[ppadder.scala 65:19]
  assign Black_21_io_i_pk = PG_13_io_s; // @[ppadder.scala 64:19]
  assign Black_21_io_i_gk = PG_13_io_co; // @[ppadder.scala 63:19]
  assign Black_22_io_i_pj = Black_21_io_o_p; // @[ppadder.scala 66:19]
  assign Black_22_io_i_gj = Black_21_io_o_g; // @[ppadder.scala 65:19]
  assign Black_22_io_i_pk = PG_14_io_s; // @[ppadder.scala 64:19]
  assign Black_22_io_i_gk = PG_14_io_co; // @[ppadder.scala 63:19]
  assign Black_23_io_i_pj = Black_22_io_o_p; // @[ppadder.scala 66:19]
  assign Black_23_io_i_gj = Black_22_io_o_g; // @[ppadder.scala 65:19]
  assign Black_23_io_i_pk = PG_15_io_s; // @[ppadder.scala 64:19]
  assign Black_23_io_i_gk = PG_15_io_co; // @[ppadder.scala 63:19]
  assign Black_24_io_i_pj = Black_23_io_o_p; // @[ppadder.scala 66:19]
  assign Black_24_io_i_gj = Black_23_io_o_g; // @[ppadder.scala 65:19]
  assign Black_24_io_i_pk = PG_16_io_s; // @[ppadder.scala 64:19]
  assign Black_24_io_i_gk = PG_16_io_co; // @[ppadder.scala 63:19]
  assign Black_25_io_i_pj = PG_10_io_s; // @[ppadder.scala 66:19]
  assign Black_25_io_i_gj = PG_10_io_co; // @[ppadder.scala 65:19]
  assign Black_25_io_i_pk = PG_11_io_s; // @[ppadder.scala 64:19]
  assign Black_25_io_i_gk = PG_11_io_co; // @[ppadder.scala 63:19]
  assign Black_26_io_i_pj = PG_7_io_s; // @[ppadder.scala 66:19]
  assign Black_26_io_i_gj = PG_7_io_co; // @[ppadder.scala 65:19]
  assign Black_26_io_i_pk = PG_8_io_s; // @[ppadder.scala 64:19]
  assign Black_26_io_i_gk = PG_8_io_co; // @[ppadder.scala 63:19]
  assign Black_27_io_i_pj = Black_26_io_o_p; // @[ppadder.scala 66:19]
  assign Black_27_io_i_gj = Black_26_io_o_g; // @[ppadder.scala 65:19]
  assign Black_27_io_i_pk = PG_9_io_s; // @[ppadder.scala 64:19]
  assign Black_27_io_i_gk = PG_9_io_co; // @[ppadder.scala 63:19]
  assign Black_28_io_i_pj = Black_27_io_o_p; // @[ppadder.scala 66:19]
  assign Black_28_io_i_gj = Black_27_io_o_g; // @[ppadder.scala 65:19]
  assign Black_28_io_i_pk = Black_25_io_o_p; // @[ppadder.scala 64:19]
  assign Black_28_io_i_gk = Black_25_io_o_g; // @[ppadder.scala 63:19]
  assign Black_29_io_i_pj = PG_5_io_s; // @[ppadder.scala 66:19]
  assign Black_29_io_i_gj = PG_5_io_co; // @[ppadder.scala 65:19]
  assign Black_29_io_i_pk = PG_6_io_s; // @[ppadder.scala 64:19]
  assign Black_29_io_i_gk = PG_6_io_co; // @[ppadder.scala 63:19]
  assign Black_30_io_i_pj = PG_4_io_s; // @[ppadder.scala 66:19]
  assign Black_30_io_i_gj = PG_4_io_co; // @[ppadder.scala 65:19]
  assign Black_30_io_i_pk = Black_29_io_o_p; // @[ppadder.scala 64:19]
  assign Black_30_io_i_gk = Black_29_io_o_g; // @[ppadder.scala 63:19]
  assign Black_31_io_i_pj = PG_2_io_s; // @[ppadder.scala 66:19]
  assign Black_31_io_i_gj = PG_2_io_co; // @[ppadder.scala 65:19]
  assign Black_31_io_i_pk = PG_3_io_s; // @[ppadder.scala 64:19]
  assign Black_31_io_i_gk = PG_3_io_co; // @[ppadder.scala 63:19]
  assign Black_32_io_i_pj = PG_io_s; // @[ppadder.scala 66:19]
  assign Black_32_io_i_gj = PG_io_co; // @[ppadder.scala 65:19]
  assign Black_32_io_i_pk = PG_1_io_s; // @[ppadder.scala 64:19]
  assign Black_32_io_i_gk = PG_1_io_co; // @[ppadder.scala 63:19]
  assign Black_33_io_i_pj = Black_32_io_o_p; // @[ppadder.scala 66:19]
  assign Black_33_io_i_gj = Black_32_io_o_g; // @[ppadder.scala 65:19]
  assign Black_33_io_i_pk = Black_31_io_o_p; // @[ppadder.scala 64:19]
  assign Black_33_io_i_gk = Black_31_io_o_g; // @[ppadder.scala 63:19]
  assign Black_34_io_i_pj = Black_33_io_o_p; // @[ppadder.scala 66:19]
  assign Black_34_io_i_gj = Black_33_io_o_g; // @[ppadder.scala 65:19]
  assign Black_34_io_i_pk = Black_30_io_o_p; // @[ppadder.scala 64:19]
  assign Black_34_io_i_gk = Black_30_io_o_g; // @[ppadder.scala 63:19]
  assign Black_35_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_35_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_35_io_i_pk = Black_28_io_o_p; // @[ppadder.scala 64:19]
  assign Black_35_io_i_gk = Black_28_io_o_g; // @[ppadder.scala 63:19]
  assign Black_36_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_36_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_36_io_i_pk = Black_24_io_o_p; // @[ppadder.scala 64:19]
  assign Black_36_io_i_gk = Black_24_io_o_g; // @[ppadder.scala 63:19]
  assign Black_37_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_37_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_37_io_i_pk = Black_12_io_o_p; // @[ppadder.scala 64:19]
  assign Black_37_io_i_gk = Black_12_io_o_g; // @[ppadder.scala 63:19]
  assign Black_38_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_38_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_38_io_i_pk = Black_13_io_o_p; // @[ppadder.scala 64:19]
  assign Black_38_io_i_gk = Black_13_io_o_g; // @[ppadder.scala 63:19]
  assign Black_39_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_39_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_39_io_i_pk = Black_14_io_o_p; // @[ppadder.scala 64:19]
  assign Black_39_io_i_gk = Black_14_io_o_g; // @[ppadder.scala 63:19]
  assign Black_40_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_40_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_40_io_i_pk = Black_15_io_o_p; // @[ppadder.scala 64:19]
  assign Black_40_io_i_gk = Black_15_io_o_g; // @[ppadder.scala 63:19]
  assign Black_41_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_41_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_41_io_i_pk = Black_16_io_o_p; // @[ppadder.scala 64:19]
  assign Black_41_io_i_gk = Black_16_io_o_g; // @[ppadder.scala 63:19]
  assign Black_42_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_42_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_42_io_i_pk = Black_11_io_o_p; // @[ppadder.scala 64:19]
  assign Black_42_io_i_gk = Black_11_io_o_g; // @[ppadder.scala 63:19]
  assign Black_43_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_43_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_43_io_i_pk = Black_17_io_o_p; // @[ppadder.scala 64:19]
  assign Black_43_io_i_gk = Black_17_io_o_g; // @[ppadder.scala 63:19]
  assign Black_44_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_44_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_44_io_i_pk = Black_18_io_o_p; // @[ppadder.scala 64:19]
  assign Black_44_io_i_gk = Black_18_io_o_g; // @[ppadder.scala 63:19]
  assign Black_45_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_45_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_45_io_i_pk = Black_19_io_o_p; // @[ppadder.scala 64:19]
  assign Black_45_io_i_gk = Black_19_io_o_g; // @[ppadder.scala 63:19]
  assign Black_46_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_46_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_46_io_i_pk = Black_10_io_o_p; // @[ppadder.scala 64:19]
  assign Black_46_io_i_gk = Black_10_io_o_g; // @[ppadder.scala 63:19]
  assign Black_47_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_47_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_47_io_i_pk = Black_20_io_o_p; // @[ppadder.scala 64:19]
  assign Black_47_io_i_gk = Black_20_io_o_g; // @[ppadder.scala 63:19]
  assign Black_48_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_48_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_48_io_i_pk = Black_9_io_o_p; // @[ppadder.scala 64:19]
  assign Black_48_io_i_gk = Black_9_io_o_g; // @[ppadder.scala 63:19]
  assign Black_49_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_49_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_49_io_i_pk = Black_8_io_o_p; // @[ppadder.scala 64:19]
  assign Black_49_io_i_gk = Black_8_io_o_g; // @[ppadder.scala 63:19]
  assign Black_50_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_50_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_50_io_i_pk = PG_17_io_s; // @[ppadder.scala 64:19]
  assign Black_50_io_i_gk = PG_17_io_co; // @[ppadder.scala 63:19]
  assign Black_51_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_51_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_51_io_i_pk = Black_23_io_o_p; // @[ppadder.scala 64:19]
  assign Black_51_io_i_gk = Black_23_io_o_g; // @[ppadder.scala 63:19]
  assign Black_52_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_52_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_52_io_i_pk = Black_22_io_o_p; // @[ppadder.scala 64:19]
  assign Black_52_io_i_gk = Black_22_io_o_g; // @[ppadder.scala 63:19]
  assign Black_53_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_53_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_53_io_i_pk = Black_21_io_o_p; // @[ppadder.scala 64:19]
  assign Black_53_io_i_gk = Black_21_io_o_g; // @[ppadder.scala 63:19]
  assign Black_54_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_54_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_54_io_i_pk = PG_12_io_s; // @[ppadder.scala 64:19]
  assign Black_54_io_i_gk = PG_12_io_co; // @[ppadder.scala 63:19]
  assign Black_55_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_55_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_55_io_i_pk = Black_27_io_o_p; // @[ppadder.scala 64:19]
  assign Black_55_io_i_gk = Black_27_io_o_g; // @[ppadder.scala 63:19]
  assign Black_56_io_i_pj = Black_55_io_o_p; // @[ppadder.scala 66:19]
  assign Black_56_io_i_gj = Black_55_io_o_g; // @[ppadder.scala 65:19]
  assign Black_56_io_i_pk = PG_10_io_s; // @[ppadder.scala 64:19]
  assign Black_56_io_i_gk = PG_10_io_co; // @[ppadder.scala 63:19]
  assign Black_57_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_57_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_57_io_i_pk = Black_26_io_o_p; // @[ppadder.scala 64:19]
  assign Black_57_io_i_gk = Black_26_io_o_g; // @[ppadder.scala 63:19]
  assign Black_58_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_58_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_58_io_i_pk = PG_7_io_s; // @[ppadder.scala 64:19]
  assign Black_58_io_i_gk = PG_7_io_co; // @[ppadder.scala 63:19]
  assign Black_59_io_i_pj = Black_33_io_o_p; // @[ppadder.scala 66:19]
  assign Black_59_io_i_gj = Black_33_io_o_g; // @[ppadder.scala 65:19]
  assign Black_59_io_i_pk = PG_4_io_s; // @[ppadder.scala 64:19]
  assign Black_59_io_i_gk = PG_4_io_co; // @[ppadder.scala 63:19]
  assign Black_60_io_i_pj = Black_59_io_o_p; // @[ppadder.scala 66:19]
  assign Black_60_io_i_gj = Black_59_io_o_g; // @[ppadder.scala 65:19]
  assign Black_60_io_i_pk = PG_5_io_s; // @[ppadder.scala 64:19]
  assign Black_60_io_i_gk = PG_5_io_co; // @[ppadder.scala 63:19]
  assign Black_61_io_i_pj = Black_32_io_o_p; // @[ppadder.scala 66:19]
  assign Black_61_io_i_gj = Black_32_io_o_g; // @[ppadder.scala 65:19]
  assign Black_61_io_i_pk = PG_2_io_s; // @[ppadder.scala 64:19]
  assign Black_61_io_i_gk = PG_2_io_co; // @[ppadder.scala 63:19]
  assign Black_62_io_i_pj = Black_37_io_o_p; // @[ppadder.scala 66:19]
  assign Black_62_io_i_gj = Black_37_io_o_g; // @[ppadder.scala 65:19]
  assign Black_62_io_i_pk = PG_31_io_s; // @[ppadder.scala 64:19]
  assign Black_62_io_i_gk = PG_31_io_co; // @[ppadder.scala 63:19]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_66) begin
          $fwrite(32'h80000002,"res(0) = %d\n",res_0); // @[ppadder.scala 77:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MACd(
  input         clock,
  input         reset,
  input  [15:0] io_multiplicand_0,
  input  [15:0] io_multiplicand_1,
  input  [15:0] io_multiplier_0,
  input  [15:0] io_multiplier_1,
  input  [31:0] io_addend,
  output [31:0] io_outs
);
  wire [15:0] pp_0_io_multiplicand; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_multiplier; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_0; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_1; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_2; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_3; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_4; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_5; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_6; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_7; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_8; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_9; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_10; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_11; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_12; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_13; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_14; // @[systolic.scala 31:48]
  wire [15:0] pp_0_io_outs_15; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_multiplicand; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_multiplier; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_0; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_1; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_2; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_3; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_4; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_5; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_6; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_7; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_8; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_9; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_10; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_11; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_12; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_13; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_14; // @[systolic.scala 31:48]
  wire [15:0] pp_1_io_outs_15; // @[systolic.scala 31:48]
  wire [15:0] wt_io_pp_0; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_1; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_2; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_3; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_4; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_5; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_6; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_7; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_8; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_9; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_10; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_11; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_12; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_13; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_14; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_15; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_16; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_17; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_18; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_19; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_20; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_21; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_22; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_23; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_24; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_25; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_26; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_27; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_28; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_29; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_30; // @[systolic.scala 37:18]
  wire [15:0] wt_io_pp_31; // @[systolic.scala 37:18]
  wire [31:0] wt_io_augend; // @[systolic.scala 37:18]
  wire [31:0] wt_io_addend; // @[systolic.scala 37:18]
  wire  ppa1_clock; // @[systolic.scala 40:20]
  wire  ppa1_reset; // @[systolic.scala 40:20]
  wire [31:0] ppa1_io_augend; // @[systolic.scala 40:20]
  wire [31:0] ppa1_io_addend; // @[systolic.scala 40:20]
  wire [31:0] ppa1_io_outs; // @[systolic.scala 40:20]
  wire  ppa2_clock; // @[systolic.scala 44:20]
  wire  ppa2_reset; // @[systolic.scala 44:20]
  wire [31:0] ppa2_io_augend; // @[systolic.scala 44:20]
  wire [31:0] ppa2_io_addend; // @[systolic.scala 44:20]
  wire [31:0] ppa2_io_outs; // @[systolic.scala 44:20]
  PartialProd pp_0 ( // @[systolic.scala 31:48]
    .io_multiplicand(pp_0_io_multiplicand),
    .io_multiplier(pp_0_io_multiplier),
    .io_outs_0(pp_0_io_outs_0),
    .io_outs_1(pp_0_io_outs_1),
    .io_outs_2(pp_0_io_outs_2),
    .io_outs_3(pp_0_io_outs_3),
    .io_outs_4(pp_0_io_outs_4),
    .io_outs_5(pp_0_io_outs_5),
    .io_outs_6(pp_0_io_outs_6),
    .io_outs_7(pp_0_io_outs_7),
    .io_outs_8(pp_0_io_outs_8),
    .io_outs_9(pp_0_io_outs_9),
    .io_outs_10(pp_0_io_outs_10),
    .io_outs_11(pp_0_io_outs_11),
    .io_outs_12(pp_0_io_outs_12),
    .io_outs_13(pp_0_io_outs_13),
    .io_outs_14(pp_0_io_outs_14),
    .io_outs_15(pp_0_io_outs_15)
  );
  PartialProd pp_1 ( // @[systolic.scala 31:48]
    .io_multiplicand(pp_1_io_multiplicand),
    .io_multiplier(pp_1_io_multiplier),
    .io_outs_0(pp_1_io_outs_0),
    .io_outs_1(pp_1_io_outs_1),
    .io_outs_2(pp_1_io_outs_2),
    .io_outs_3(pp_1_io_outs_3),
    .io_outs_4(pp_1_io_outs_4),
    .io_outs_5(pp_1_io_outs_5),
    .io_outs_6(pp_1_io_outs_6),
    .io_outs_7(pp_1_io_outs_7),
    .io_outs_8(pp_1_io_outs_8),
    .io_outs_9(pp_1_io_outs_9),
    .io_outs_10(pp_1_io_outs_10),
    .io_outs_11(pp_1_io_outs_11),
    .io_outs_12(pp_1_io_outs_12),
    .io_outs_13(pp_1_io_outs_13),
    .io_outs_14(pp_1_io_outs_14),
    .io_outs_15(pp_1_io_outs_15)
  );
  Wallaced wt ( // @[systolic.scala 37:18]
    .io_pp_0(wt_io_pp_0),
    .io_pp_1(wt_io_pp_1),
    .io_pp_2(wt_io_pp_2),
    .io_pp_3(wt_io_pp_3),
    .io_pp_4(wt_io_pp_4),
    .io_pp_5(wt_io_pp_5),
    .io_pp_6(wt_io_pp_6),
    .io_pp_7(wt_io_pp_7),
    .io_pp_8(wt_io_pp_8),
    .io_pp_9(wt_io_pp_9),
    .io_pp_10(wt_io_pp_10),
    .io_pp_11(wt_io_pp_11),
    .io_pp_12(wt_io_pp_12),
    .io_pp_13(wt_io_pp_13),
    .io_pp_14(wt_io_pp_14),
    .io_pp_15(wt_io_pp_15),
    .io_pp_16(wt_io_pp_16),
    .io_pp_17(wt_io_pp_17),
    .io_pp_18(wt_io_pp_18),
    .io_pp_19(wt_io_pp_19),
    .io_pp_20(wt_io_pp_20),
    .io_pp_21(wt_io_pp_21),
    .io_pp_22(wt_io_pp_22),
    .io_pp_23(wt_io_pp_23),
    .io_pp_24(wt_io_pp_24),
    .io_pp_25(wt_io_pp_25),
    .io_pp_26(wt_io_pp_26),
    .io_pp_27(wt_io_pp_27),
    .io_pp_28(wt_io_pp_28),
    .io_pp_29(wt_io_pp_29),
    .io_pp_30(wt_io_pp_30),
    .io_pp_31(wt_io_pp_31),
    .io_augend(wt_io_augend),
    .io_addend(wt_io_addend)
  );
  PPAdder ppa1 ( // @[systolic.scala 40:20]
    .clock(ppa1_clock),
    .reset(ppa1_reset),
    .io_augend(ppa1_io_augend),
    .io_addend(ppa1_io_addend),
    .io_outs(ppa1_io_outs)
  );
  PPAdder ppa2 ( // @[systolic.scala 44:20]
    .clock(ppa2_clock),
    .reset(ppa2_reset),
    .io_augend(ppa2_io_augend),
    .io_addend(ppa2_io_addend),
    .io_outs(ppa2_io_outs)
  );
  assign io_outs = ppa2_io_outs; // @[systolic.scala 48:11]
  assign pp_0_io_multiplicand = io_multiplicand_0; // @[systolic.scala 33:27]
  assign pp_0_io_multiplier = io_multiplier_0; // @[systolic.scala 34:25]
  assign pp_1_io_multiplicand = io_multiplicand_1; // @[systolic.scala 33:27]
  assign pp_1_io_multiplier = io_multiplier_1; // @[systolic.scala 34:25]
  assign wt_io_pp_0 = pp_0_io_outs_0; // @[systolic.scala 39:12]
  assign wt_io_pp_1 = pp_0_io_outs_1; // @[systolic.scala 39:12]
  assign wt_io_pp_2 = pp_0_io_outs_2; // @[systolic.scala 39:12]
  assign wt_io_pp_3 = pp_0_io_outs_3; // @[systolic.scala 39:12]
  assign wt_io_pp_4 = pp_0_io_outs_4; // @[systolic.scala 39:12]
  assign wt_io_pp_5 = pp_0_io_outs_5; // @[systolic.scala 39:12]
  assign wt_io_pp_6 = pp_0_io_outs_6; // @[systolic.scala 39:12]
  assign wt_io_pp_7 = pp_0_io_outs_7; // @[systolic.scala 39:12]
  assign wt_io_pp_8 = pp_0_io_outs_8; // @[systolic.scala 39:12]
  assign wt_io_pp_9 = pp_0_io_outs_9; // @[systolic.scala 39:12]
  assign wt_io_pp_10 = pp_0_io_outs_10; // @[systolic.scala 39:12]
  assign wt_io_pp_11 = pp_0_io_outs_11; // @[systolic.scala 39:12]
  assign wt_io_pp_12 = pp_0_io_outs_12; // @[systolic.scala 39:12]
  assign wt_io_pp_13 = pp_0_io_outs_13; // @[systolic.scala 39:12]
  assign wt_io_pp_14 = pp_0_io_outs_14; // @[systolic.scala 39:12]
  assign wt_io_pp_15 = pp_0_io_outs_15; // @[systolic.scala 39:12]
  assign wt_io_pp_16 = pp_1_io_outs_0; // @[systolic.scala 39:12]
  assign wt_io_pp_17 = pp_1_io_outs_1; // @[systolic.scala 39:12]
  assign wt_io_pp_18 = pp_1_io_outs_2; // @[systolic.scala 39:12]
  assign wt_io_pp_19 = pp_1_io_outs_3; // @[systolic.scala 39:12]
  assign wt_io_pp_20 = pp_1_io_outs_4; // @[systolic.scala 39:12]
  assign wt_io_pp_21 = pp_1_io_outs_5; // @[systolic.scala 39:12]
  assign wt_io_pp_22 = pp_1_io_outs_6; // @[systolic.scala 39:12]
  assign wt_io_pp_23 = pp_1_io_outs_7; // @[systolic.scala 39:12]
  assign wt_io_pp_24 = pp_1_io_outs_8; // @[systolic.scala 39:12]
  assign wt_io_pp_25 = pp_1_io_outs_9; // @[systolic.scala 39:12]
  assign wt_io_pp_26 = pp_1_io_outs_10; // @[systolic.scala 39:12]
  assign wt_io_pp_27 = pp_1_io_outs_11; // @[systolic.scala 39:12]
  assign wt_io_pp_28 = pp_1_io_outs_12; // @[systolic.scala 39:12]
  assign wt_io_pp_29 = pp_1_io_outs_13; // @[systolic.scala 39:12]
  assign wt_io_pp_30 = pp_1_io_outs_14; // @[systolic.scala 39:12]
  assign wt_io_pp_31 = pp_1_io_outs_15; // @[systolic.scala 39:12]
  assign ppa1_clock = clock;
  assign ppa1_reset = reset;
  assign ppa1_io_augend = wt_io_augend; // @[systolic.scala 41:18]
  assign ppa1_io_addend = wt_io_addend; // @[systolic.scala 42:18]
  assign ppa2_clock = clock;
  assign ppa2_reset = reset;
  assign ppa2_io_augend = ppa1_io_outs; // @[systolic.scala 45:18]
  assign ppa2_io_addend = io_addend; // @[systolic.scala 46:18]
endmodule
