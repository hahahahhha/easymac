module PartialProd(
  input  [15:0] io_multiplicand,
  input  [15:0] io_multiplier,
  output [15:0] io_outs_0,
  output [15:0] io_outs_1,
  output [15:0] io_outs_2,
  output [15:0] io_outs_3,
  output [15:0] io_outs_4,
  output [15:0] io_outs_5,
  output [15:0] io_outs_6,
  output [15:0] io_outs_7,
  output [15:0] io_outs_8,
  output [15:0] io_outs_9,
  output [15:0] io_outs_10,
  output [15:0] io_outs_11,
  output [15:0] io_outs_12,
  output [15:0] io_outs_13,
  output [15:0] io_outs_14,
  output [15:0] io_outs_15
);
  wire  _T_18 = io_multiplicand[0] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_21 = io_multiplicand[1] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_24 = io_multiplicand[2] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_27 = io_multiplicand[3] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_30 = io_multiplicand[4] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_33 = io_multiplicand[5] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_36 = io_multiplicand[6] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_39 = io_multiplicand[7] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_42 = io_multiplicand[8] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_45 = io_multiplicand[9] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_48 = io_multiplicand[10] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_51 = io_multiplicand[11] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_54 = io_multiplicand[12] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_57 = io_multiplicand[13] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_60 = io_multiplicand[14] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire  _T_63 = io_multiplicand[15] & io_multiplier[0]; // @[partialprod.scala 16:36]
  wire [9:0] _T_72 = {_T_63,_T_60,_T_57,_T_54,_T_51,_T_48,_T_45,_T_42,_T_39,_T_36}; // @[Cat.scala 29:58]
  wire [14:0] _T_77 = {_T_72,_T_33,_T_30,_T_27,_T_24,_T_21}; // @[Cat.scala 29:58]
  wire  _T_97 = io_multiplicand[0] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_100 = io_multiplicand[1] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_103 = io_multiplicand[2] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_106 = io_multiplicand[3] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_109 = io_multiplicand[4] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_112 = io_multiplicand[5] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_115 = io_multiplicand[6] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_118 = io_multiplicand[7] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_121 = io_multiplicand[8] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_124 = io_multiplicand[9] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_127 = io_multiplicand[10] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_130 = io_multiplicand[11] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_133 = io_multiplicand[12] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_136 = io_multiplicand[13] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_139 = io_multiplicand[14] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire  _T_142 = io_multiplicand[15] & io_multiplier[1]; // @[partialprod.scala 16:36]
  wire [9:0] _T_151 = {_T_142,_T_139,_T_136,_T_133,_T_130,_T_127,_T_124,_T_121,_T_118,_T_115}; // @[Cat.scala 29:58]
  wire [14:0] _T_156 = {_T_151,_T_112,_T_109,_T_106,_T_103,_T_100}; // @[Cat.scala 29:58]
  wire  _T_176 = io_multiplicand[0] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_179 = io_multiplicand[1] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_182 = io_multiplicand[2] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_185 = io_multiplicand[3] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_188 = io_multiplicand[4] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_191 = io_multiplicand[5] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_194 = io_multiplicand[6] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_197 = io_multiplicand[7] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_200 = io_multiplicand[8] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_203 = io_multiplicand[9] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_206 = io_multiplicand[10] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_209 = io_multiplicand[11] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_212 = io_multiplicand[12] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_215 = io_multiplicand[13] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_218 = io_multiplicand[14] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire  _T_221 = io_multiplicand[15] & io_multiplier[2]; // @[partialprod.scala 16:36]
  wire [9:0] _T_230 = {_T_221,_T_218,_T_215,_T_212,_T_209,_T_206,_T_203,_T_200,_T_197,_T_194}; // @[Cat.scala 29:58]
  wire [14:0] _T_235 = {_T_230,_T_191,_T_188,_T_185,_T_182,_T_179}; // @[Cat.scala 29:58]
  wire  _T_255 = io_multiplicand[0] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_258 = io_multiplicand[1] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_261 = io_multiplicand[2] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_264 = io_multiplicand[3] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_267 = io_multiplicand[4] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_270 = io_multiplicand[5] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_273 = io_multiplicand[6] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_276 = io_multiplicand[7] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_279 = io_multiplicand[8] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_282 = io_multiplicand[9] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_285 = io_multiplicand[10] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_288 = io_multiplicand[11] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_291 = io_multiplicand[12] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_294 = io_multiplicand[13] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_297 = io_multiplicand[14] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire  _T_300 = io_multiplicand[15] & io_multiplier[3]; // @[partialprod.scala 16:36]
  wire [9:0] _T_309 = {_T_300,_T_297,_T_294,_T_291,_T_288,_T_285,_T_282,_T_279,_T_276,_T_273}; // @[Cat.scala 29:58]
  wire [14:0] _T_314 = {_T_309,_T_270,_T_267,_T_264,_T_261,_T_258}; // @[Cat.scala 29:58]
  wire  _T_334 = io_multiplicand[0] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_337 = io_multiplicand[1] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_340 = io_multiplicand[2] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_343 = io_multiplicand[3] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_346 = io_multiplicand[4] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_349 = io_multiplicand[5] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_352 = io_multiplicand[6] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_355 = io_multiplicand[7] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_358 = io_multiplicand[8] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_361 = io_multiplicand[9] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_364 = io_multiplicand[10] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_367 = io_multiplicand[11] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_370 = io_multiplicand[12] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_373 = io_multiplicand[13] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_376 = io_multiplicand[14] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire  _T_379 = io_multiplicand[15] & io_multiplier[4]; // @[partialprod.scala 16:36]
  wire [9:0] _T_388 = {_T_379,_T_376,_T_373,_T_370,_T_367,_T_364,_T_361,_T_358,_T_355,_T_352}; // @[Cat.scala 29:58]
  wire [14:0] _T_393 = {_T_388,_T_349,_T_346,_T_343,_T_340,_T_337}; // @[Cat.scala 29:58]
  wire  _T_413 = io_multiplicand[0] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_416 = io_multiplicand[1] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_419 = io_multiplicand[2] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_422 = io_multiplicand[3] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_425 = io_multiplicand[4] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_428 = io_multiplicand[5] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_431 = io_multiplicand[6] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_434 = io_multiplicand[7] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_437 = io_multiplicand[8] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_440 = io_multiplicand[9] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_443 = io_multiplicand[10] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_446 = io_multiplicand[11] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_449 = io_multiplicand[12] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_452 = io_multiplicand[13] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_455 = io_multiplicand[14] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire  _T_458 = io_multiplicand[15] & io_multiplier[5]; // @[partialprod.scala 16:36]
  wire [9:0] _T_467 = {_T_458,_T_455,_T_452,_T_449,_T_446,_T_443,_T_440,_T_437,_T_434,_T_431}; // @[Cat.scala 29:58]
  wire [14:0] _T_472 = {_T_467,_T_428,_T_425,_T_422,_T_419,_T_416}; // @[Cat.scala 29:58]
  wire  _T_492 = io_multiplicand[0] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_495 = io_multiplicand[1] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_498 = io_multiplicand[2] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_501 = io_multiplicand[3] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_504 = io_multiplicand[4] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_507 = io_multiplicand[5] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_510 = io_multiplicand[6] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_513 = io_multiplicand[7] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_516 = io_multiplicand[8] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_519 = io_multiplicand[9] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_522 = io_multiplicand[10] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_525 = io_multiplicand[11] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_528 = io_multiplicand[12] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_531 = io_multiplicand[13] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_534 = io_multiplicand[14] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire  _T_537 = io_multiplicand[15] & io_multiplier[6]; // @[partialprod.scala 16:36]
  wire [9:0] _T_546 = {_T_537,_T_534,_T_531,_T_528,_T_525,_T_522,_T_519,_T_516,_T_513,_T_510}; // @[Cat.scala 29:58]
  wire [14:0] _T_551 = {_T_546,_T_507,_T_504,_T_501,_T_498,_T_495}; // @[Cat.scala 29:58]
  wire  _T_571 = io_multiplicand[0] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_574 = io_multiplicand[1] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_577 = io_multiplicand[2] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_580 = io_multiplicand[3] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_583 = io_multiplicand[4] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_586 = io_multiplicand[5] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_589 = io_multiplicand[6] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_592 = io_multiplicand[7] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_595 = io_multiplicand[8] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_598 = io_multiplicand[9] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_601 = io_multiplicand[10] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_604 = io_multiplicand[11] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_607 = io_multiplicand[12] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_610 = io_multiplicand[13] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_613 = io_multiplicand[14] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire  _T_616 = io_multiplicand[15] & io_multiplier[7]; // @[partialprod.scala 16:36]
  wire [9:0] _T_625 = {_T_616,_T_613,_T_610,_T_607,_T_604,_T_601,_T_598,_T_595,_T_592,_T_589}; // @[Cat.scala 29:58]
  wire [14:0] _T_630 = {_T_625,_T_586,_T_583,_T_580,_T_577,_T_574}; // @[Cat.scala 29:58]
  wire  _T_650 = io_multiplicand[0] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_653 = io_multiplicand[1] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_656 = io_multiplicand[2] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_659 = io_multiplicand[3] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_662 = io_multiplicand[4] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_665 = io_multiplicand[5] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_668 = io_multiplicand[6] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_671 = io_multiplicand[7] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_674 = io_multiplicand[8] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_677 = io_multiplicand[9] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_680 = io_multiplicand[10] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_683 = io_multiplicand[11] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_686 = io_multiplicand[12] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_689 = io_multiplicand[13] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_692 = io_multiplicand[14] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire  _T_695 = io_multiplicand[15] & io_multiplier[8]; // @[partialprod.scala 16:36]
  wire [9:0] _T_704 = {_T_695,_T_692,_T_689,_T_686,_T_683,_T_680,_T_677,_T_674,_T_671,_T_668}; // @[Cat.scala 29:58]
  wire [14:0] _T_709 = {_T_704,_T_665,_T_662,_T_659,_T_656,_T_653}; // @[Cat.scala 29:58]
  wire  _T_729 = io_multiplicand[0] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_732 = io_multiplicand[1] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_735 = io_multiplicand[2] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_738 = io_multiplicand[3] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_741 = io_multiplicand[4] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_744 = io_multiplicand[5] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_747 = io_multiplicand[6] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_750 = io_multiplicand[7] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_753 = io_multiplicand[8] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_756 = io_multiplicand[9] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_759 = io_multiplicand[10] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_762 = io_multiplicand[11] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_765 = io_multiplicand[12] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_768 = io_multiplicand[13] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_771 = io_multiplicand[14] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire  _T_774 = io_multiplicand[15] & io_multiplier[9]; // @[partialprod.scala 16:36]
  wire [9:0] _T_783 = {_T_774,_T_771,_T_768,_T_765,_T_762,_T_759,_T_756,_T_753,_T_750,_T_747}; // @[Cat.scala 29:58]
  wire [14:0] _T_788 = {_T_783,_T_744,_T_741,_T_738,_T_735,_T_732}; // @[Cat.scala 29:58]
  wire  _T_808 = io_multiplicand[0] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_811 = io_multiplicand[1] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_814 = io_multiplicand[2] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_817 = io_multiplicand[3] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_820 = io_multiplicand[4] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_823 = io_multiplicand[5] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_826 = io_multiplicand[6] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_829 = io_multiplicand[7] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_832 = io_multiplicand[8] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_835 = io_multiplicand[9] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_838 = io_multiplicand[10] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_841 = io_multiplicand[11] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_844 = io_multiplicand[12] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_847 = io_multiplicand[13] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_850 = io_multiplicand[14] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire  _T_853 = io_multiplicand[15] & io_multiplier[10]; // @[partialprod.scala 16:36]
  wire [9:0] _T_862 = {_T_853,_T_850,_T_847,_T_844,_T_841,_T_838,_T_835,_T_832,_T_829,_T_826}; // @[Cat.scala 29:58]
  wire [14:0] _T_867 = {_T_862,_T_823,_T_820,_T_817,_T_814,_T_811}; // @[Cat.scala 29:58]
  wire  _T_887 = io_multiplicand[0] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_890 = io_multiplicand[1] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_893 = io_multiplicand[2] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_896 = io_multiplicand[3] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_899 = io_multiplicand[4] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_902 = io_multiplicand[5] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_905 = io_multiplicand[6] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_908 = io_multiplicand[7] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_911 = io_multiplicand[8] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_914 = io_multiplicand[9] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_917 = io_multiplicand[10] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_920 = io_multiplicand[11] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_923 = io_multiplicand[12] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_926 = io_multiplicand[13] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_929 = io_multiplicand[14] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire  _T_932 = io_multiplicand[15] & io_multiplier[11]; // @[partialprod.scala 16:36]
  wire [9:0] _T_941 = {_T_932,_T_929,_T_926,_T_923,_T_920,_T_917,_T_914,_T_911,_T_908,_T_905}; // @[Cat.scala 29:58]
  wire [14:0] _T_946 = {_T_941,_T_902,_T_899,_T_896,_T_893,_T_890}; // @[Cat.scala 29:58]
  wire  _T_966 = io_multiplicand[0] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_969 = io_multiplicand[1] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_972 = io_multiplicand[2] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_975 = io_multiplicand[3] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_978 = io_multiplicand[4] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_981 = io_multiplicand[5] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_984 = io_multiplicand[6] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_987 = io_multiplicand[7] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_990 = io_multiplicand[8] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_993 = io_multiplicand[9] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_996 = io_multiplicand[10] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_999 = io_multiplicand[11] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1002 = io_multiplicand[12] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1005 = io_multiplicand[13] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1008 = io_multiplicand[14] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire  _T_1011 = io_multiplicand[15] & io_multiplier[12]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1020 = {_T_1011,_T_1008,_T_1005,_T_1002,_T_999,_T_996,_T_993,_T_990,_T_987,_T_984}; // @[Cat.scala 29:58]
  wire [14:0] _T_1025 = {_T_1020,_T_981,_T_978,_T_975,_T_972,_T_969}; // @[Cat.scala 29:58]
  wire  _T_1045 = io_multiplicand[0] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1048 = io_multiplicand[1] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1051 = io_multiplicand[2] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1054 = io_multiplicand[3] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1057 = io_multiplicand[4] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1060 = io_multiplicand[5] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1063 = io_multiplicand[6] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1066 = io_multiplicand[7] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1069 = io_multiplicand[8] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1072 = io_multiplicand[9] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1075 = io_multiplicand[10] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1078 = io_multiplicand[11] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1081 = io_multiplicand[12] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1084 = io_multiplicand[13] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1087 = io_multiplicand[14] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire  _T_1090 = io_multiplicand[15] & io_multiplier[13]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1099 = {_T_1090,_T_1087,_T_1084,_T_1081,_T_1078,_T_1075,_T_1072,_T_1069,_T_1066,_T_1063}; // @[Cat.scala 29:58]
  wire [14:0] _T_1104 = {_T_1099,_T_1060,_T_1057,_T_1054,_T_1051,_T_1048}; // @[Cat.scala 29:58]
  wire  _T_1124 = io_multiplicand[0] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1127 = io_multiplicand[1] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1130 = io_multiplicand[2] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1133 = io_multiplicand[3] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1136 = io_multiplicand[4] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1139 = io_multiplicand[5] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1142 = io_multiplicand[6] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1145 = io_multiplicand[7] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1148 = io_multiplicand[8] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1151 = io_multiplicand[9] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1154 = io_multiplicand[10] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1157 = io_multiplicand[11] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1160 = io_multiplicand[12] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1163 = io_multiplicand[13] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1166 = io_multiplicand[14] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire  _T_1169 = io_multiplicand[15] & io_multiplier[14]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1178 = {_T_1169,_T_1166,_T_1163,_T_1160,_T_1157,_T_1154,_T_1151,_T_1148,_T_1145,_T_1142}; // @[Cat.scala 29:58]
  wire [14:0] _T_1183 = {_T_1178,_T_1139,_T_1136,_T_1133,_T_1130,_T_1127}; // @[Cat.scala 29:58]
  wire  _T_1203 = io_multiplicand[0] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1206 = io_multiplicand[1] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1209 = io_multiplicand[2] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1212 = io_multiplicand[3] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1215 = io_multiplicand[4] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1218 = io_multiplicand[5] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1221 = io_multiplicand[6] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1224 = io_multiplicand[7] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1227 = io_multiplicand[8] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1230 = io_multiplicand[9] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1233 = io_multiplicand[10] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1236 = io_multiplicand[11] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1239 = io_multiplicand[12] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1242 = io_multiplicand[13] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1245 = io_multiplicand[14] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire  _T_1248 = io_multiplicand[15] & io_multiplier[15]; // @[partialprod.scala 16:36]
  wire [9:0] _T_1257 = {_T_1248,_T_1245,_T_1242,_T_1239,_T_1236,_T_1233,_T_1230,_T_1227,_T_1224,_T_1221}; // @[Cat.scala 29:58]
  wire [14:0] _T_1262 = {_T_1257,_T_1218,_T_1215,_T_1212,_T_1209,_T_1206}; // @[Cat.scala 29:58]
  assign io_outs_0 = {_T_77,_T_18}; // @[partialprod.scala 18:16]
  assign io_outs_1 = {_T_156,_T_97}; // @[partialprod.scala 18:16]
  assign io_outs_2 = {_T_235,_T_176}; // @[partialprod.scala 18:16]
  assign io_outs_3 = {_T_314,_T_255}; // @[partialprod.scala 18:16]
  assign io_outs_4 = {_T_393,_T_334}; // @[partialprod.scala 18:16]
  assign io_outs_5 = {_T_472,_T_413}; // @[partialprod.scala 18:16]
  assign io_outs_6 = {_T_551,_T_492}; // @[partialprod.scala 18:16]
  assign io_outs_7 = {_T_630,_T_571}; // @[partialprod.scala 18:16]
  assign io_outs_8 = {_T_709,_T_650}; // @[partialprod.scala 18:16]
  assign io_outs_9 = {_T_788,_T_729}; // @[partialprod.scala 18:16]
  assign io_outs_10 = {_T_867,_T_808}; // @[partialprod.scala 18:16]
  assign io_outs_11 = {_T_946,_T_887}; // @[partialprod.scala 18:16]
  assign io_outs_12 = {_T_1025,_T_966}; // @[partialprod.scala 18:16]
  assign io_outs_13 = {_T_1104,_T_1045}; // @[partialprod.scala 18:16]
  assign io_outs_14 = {_T_1183,_T_1124}; // @[partialprod.scala 18:16]
  assign io_outs_15 = {_T_1262,_T_1203}; // @[partialprod.scala 18:16]
endmodule
module FullAdder(
  input   io_a,
  input   io_b,
  input   io_ci,
  output  io_s,
  output  io_co
);
  wire  a_xor_b = io_a ^ io_b; // @[comp.scala 28:22]
  wire  a_and_b = io_a & io_b; // @[comp.scala 31:22]
  wire  a_and_cin = io_a & io_ci; // @[comp.scala 32:24]
  wire  b_and_cin = io_b & io_ci; // @[comp.scala 33:24]
  wire  _T_1 = a_and_b | b_and_cin; // @[comp.scala 34:20]
  assign io_s = a_xor_b ^ io_ci; // @[comp.scala 29:8]
  assign io_co = _T_1 | a_and_cin; // @[comp.scala 34:9]
endmodule
module HalfAdder(
  input   io_a,
  input   io_b,
  output  io_s,
  output  io_co
);
  assign io_s = io_a ^ io_b; // @[comp.scala 15:8]
  assign io_co = io_a & io_b; // @[comp.scala 16:9]
endmodule
module Wallace(
  input  [15:0] io_pp_0,
  input  [15:0] io_pp_1,
  input  [15:0] io_pp_2,
  input  [15:0] io_pp_3,
  input  [15:0] io_pp_4,
  input  [15:0] io_pp_5,
  input  [15:0] io_pp_6,
  input  [15:0] io_pp_7,
  input  [15:0] io_pp_8,
  input  [15:0] io_pp_9,
  input  [15:0] io_pp_10,
  input  [15:0] io_pp_11,
  input  [15:0] io_pp_12,
  input  [15:0] io_pp_13,
  input  [15:0] io_pp_14,
  input  [15:0] io_pp_15,
  output [31:0] io_augend,
  output [31:0] io_addend
);
  wire  FullAdder_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_1_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_1_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_1_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_1_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_1_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_2_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_2_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_2_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_2_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_2_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_3_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_3_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_3_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_3_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_3_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_4_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_4_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_4_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_4_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_4_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_5_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_5_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_5_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_5_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_5_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_6_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_6_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_6_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_6_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_6_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_7_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_7_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_7_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_7_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_7_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_8_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_8_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_8_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_8_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_8_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_9_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_9_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_9_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_9_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_9_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_10_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_10_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_10_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_10_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_10_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_11_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_11_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_11_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_11_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_11_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_12_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_12_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_12_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_12_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_12_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_13_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_13_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_13_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_13_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_13_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_14_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_14_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_14_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_14_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_14_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_15_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_15_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_15_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_15_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_15_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_16_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_16_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_16_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_16_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_16_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_17_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_17_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_17_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_17_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_17_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_18_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_18_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_18_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_18_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_18_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_19_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_19_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_19_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_19_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_19_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_20_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_20_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_20_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_20_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_20_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_21_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_21_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_21_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_21_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_21_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_22_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_22_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_22_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_22_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_22_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_23_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_23_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_23_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_23_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_23_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_24_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_24_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_24_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_24_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_24_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_25_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_25_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_25_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_25_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_25_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_26_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_26_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_26_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_26_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_26_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_27_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_27_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_27_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_27_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_27_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_28_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_28_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_28_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_28_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_28_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_29_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_29_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_29_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_29_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_29_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_30_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_30_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_30_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_30_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_30_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_31_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_31_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_31_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_31_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_31_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_32_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_32_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_32_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_32_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_32_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_33_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_33_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_33_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_33_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_33_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_34_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_34_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_34_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_34_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_34_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_35_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_35_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_35_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_35_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_35_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_36_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_36_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_36_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_36_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_36_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_37_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_37_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_37_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_37_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_37_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_38_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_38_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_38_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_38_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_38_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_39_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_39_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_39_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_39_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_39_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_40_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_40_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_40_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_40_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_40_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_41_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_41_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_41_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_41_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_41_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_42_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_42_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_42_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_42_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_42_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_43_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_43_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_43_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_43_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_43_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_44_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_44_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_44_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_44_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_44_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_45_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_45_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_45_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_45_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_45_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_46_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_46_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_46_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_46_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_46_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_47_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_47_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_47_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_47_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_47_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_48_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_48_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_48_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_48_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_48_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_49_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_49_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_49_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_49_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_49_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_50_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_50_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_50_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_50_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_50_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_51_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_51_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_51_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_51_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_51_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_52_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_52_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_52_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_52_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_52_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_53_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_53_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_53_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_53_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_53_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_54_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_54_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_54_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_54_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_54_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_55_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_55_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_55_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_55_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_55_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_56_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_56_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_56_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_56_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_56_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_57_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_57_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_57_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_57_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_57_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_58_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_58_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_58_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_58_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_58_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_59_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_59_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_59_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_59_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_59_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_60_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_60_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_60_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_60_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_60_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_61_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_61_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_61_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_61_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_61_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_62_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_62_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_62_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_62_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_62_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_63_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_63_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_63_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_63_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_63_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_64_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_64_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_64_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_64_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_64_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_65_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_65_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_65_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_65_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_65_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_66_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_66_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_66_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_66_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_66_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_67_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_67_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_67_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_67_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_67_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_68_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_68_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_68_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_68_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_68_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_69_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_69_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_69_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_69_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_69_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_70_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_70_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_70_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_70_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_70_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_71_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_71_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_71_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_71_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_71_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_72_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_72_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_72_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_72_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_72_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_73_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_73_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_73_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_73_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_73_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_74_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_74_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_74_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_74_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_74_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_75_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_75_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_75_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_75_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_75_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_76_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_76_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_76_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_76_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_76_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_77_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_77_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_77_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_77_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_77_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_78_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_78_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_78_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_78_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_78_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_79_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_79_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_79_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_79_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_79_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_80_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_80_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_80_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_80_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_80_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_81_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_81_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_81_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_81_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_81_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_82_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_82_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_82_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_82_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_82_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_83_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_83_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_83_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_83_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_83_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_84_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_84_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_84_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_84_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_84_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_85_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_85_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_85_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_85_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_85_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_86_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_86_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_86_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_86_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_86_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_87_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_87_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_87_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_87_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_87_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_88_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_88_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_88_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_88_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_88_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_89_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_89_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_89_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_89_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_89_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_90_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_90_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_90_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_90_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_90_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_91_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_91_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_91_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_91_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_91_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_92_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_92_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_92_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_92_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_92_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_93_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_93_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_93_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_93_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_93_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_94_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_94_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_94_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_94_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_94_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_95_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_95_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_95_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_95_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_95_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_96_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_96_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_96_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_96_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_96_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_97_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_97_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_97_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_97_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_97_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_98_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_98_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_98_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_98_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_98_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_99_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_99_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_99_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_99_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_99_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_100_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_100_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_100_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_100_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_100_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_101_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_101_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_101_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_101_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_101_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_102_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_102_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_102_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_102_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_102_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_103_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_103_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_103_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_103_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_103_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_104_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_104_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_104_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_104_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_104_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_105_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_105_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_105_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_105_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_105_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_106_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_106_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_106_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_106_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_106_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_107_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_107_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_107_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_107_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_107_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_108_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_108_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_108_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_108_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_108_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_109_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_109_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_109_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_109_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_109_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_110_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_110_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_110_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_110_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_110_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_111_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_111_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_111_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_111_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_111_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_112_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_112_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_112_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_112_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_112_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_113_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_113_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_113_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_113_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_113_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_114_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_114_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_114_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_114_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_114_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_115_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_115_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_115_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_115_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_115_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_116_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_116_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_116_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_116_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_116_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_117_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_117_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_117_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_117_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_117_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_118_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_118_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_118_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_118_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_118_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_119_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_119_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_119_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_119_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_119_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_120_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_120_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_120_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_120_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_120_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_121_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_121_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_121_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_121_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_121_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_122_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_122_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_122_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_122_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_122_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_123_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_123_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_123_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_123_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_123_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_124_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_124_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_124_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_124_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_124_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_125_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_125_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_125_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_125_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_125_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_126_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_126_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_126_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_126_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_126_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_127_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_127_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_127_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_127_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_127_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_128_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_128_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_128_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_128_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_128_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_129_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_129_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_129_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_129_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_129_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_130_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_130_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_130_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_130_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_130_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_131_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_131_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_131_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_131_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_131_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_132_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_132_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_132_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_132_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_132_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_133_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_133_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_133_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_133_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_133_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_134_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_134_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_134_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_134_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_134_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_135_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_135_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_135_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_135_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_135_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_136_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_136_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_136_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_136_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_136_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_137_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_137_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_137_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_137_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_137_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_138_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_138_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_138_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_138_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_138_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_139_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_139_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_139_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_139_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_139_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_140_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_140_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_140_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_140_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_140_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_141_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_141_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_141_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_141_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_141_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_142_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_142_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_142_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_142_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_142_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_143_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_143_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_143_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_143_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_143_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_144_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_144_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_144_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_144_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_144_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_145_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_145_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_145_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_145_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_145_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_146_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_146_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_146_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_146_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_146_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_147_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_147_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_147_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_147_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_147_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_148_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_148_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_148_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_148_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_148_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_149_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_149_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_149_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_149_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_149_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_150_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_150_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_150_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_150_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_150_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_151_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_151_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_151_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_151_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_151_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_152_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_152_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_152_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_152_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_152_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_153_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_153_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_153_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_153_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_153_io_co; // @[wallace.scala 63:25]
  wire  HalfAdder_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_io_co; // @[wallace.scala 54:25]
  wire  FullAdder_154_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_154_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_154_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_154_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_154_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_155_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_155_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_155_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_155_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_155_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_156_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_156_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_156_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_156_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_156_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_157_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_157_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_157_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_157_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_157_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_158_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_158_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_158_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_158_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_158_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_159_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_159_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_159_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_159_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_159_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_160_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_160_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_160_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_160_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_160_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_161_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_161_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_161_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_161_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_161_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_162_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_162_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_162_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_162_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_162_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_163_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_163_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_163_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_163_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_163_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_164_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_164_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_164_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_164_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_164_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_165_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_165_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_165_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_165_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_165_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_166_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_166_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_166_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_166_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_166_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_167_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_167_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_167_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_167_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_167_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_168_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_168_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_168_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_168_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_168_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_169_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_169_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_169_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_169_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_169_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_170_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_170_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_170_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_170_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_170_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_171_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_171_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_171_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_171_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_171_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_172_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_172_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_172_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_172_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_172_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_173_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_173_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_173_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_173_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_173_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_174_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_174_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_174_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_174_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_174_io_co; // @[wallace.scala 63:25]
  wire  HalfAdder_1_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_1_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_1_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_1_io_co; // @[wallace.scala 54:25]
  wire  FullAdder_175_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_175_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_175_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_175_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_175_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_176_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_176_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_176_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_176_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_176_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_177_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_177_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_177_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_177_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_177_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_178_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_178_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_178_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_178_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_178_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_179_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_179_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_179_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_179_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_179_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_180_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_180_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_180_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_180_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_180_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_181_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_181_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_181_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_181_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_181_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_182_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_182_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_182_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_182_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_182_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_183_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_183_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_183_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_183_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_183_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_184_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_184_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_184_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_184_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_184_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_185_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_185_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_185_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_185_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_185_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_186_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_186_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_186_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_186_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_186_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_187_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_187_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_187_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_187_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_187_io_co; // @[wallace.scala 63:25]
  wire  HalfAdder_2_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_2_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_2_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_2_io_co; // @[wallace.scala 54:25]
  wire  FullAdder_188_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_188_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_188_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_188_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_188_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_189_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_189_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_189_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_189_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_189_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_190_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_190_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_190_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_190_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_190_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_191_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_191_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_191_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_191_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_191_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_192_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_192_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_192_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_192_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_192_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_193_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_193_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_193_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_193_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_193_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_194_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_194_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_194_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_194_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_194_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_195_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_195_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_195_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_195_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_195_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_196_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_196_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_196_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_196_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_196_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_197_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_197_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_197_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_197_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_197_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_198_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_198_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_198_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_198_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_198_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_199_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_199_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_199_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_199_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_199_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_200_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_200_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_200_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_200_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_200_io_co; // @[wallace.scala 63:25]
  wire  HalfAdder_3_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_3_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_3_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_3_io_co; // @[wallace.scala 54:25]
  wire  HalfAdder_4_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_4_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_4_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_4_io_co; // @[wallace.scala 54:25]
  wire  HalfAdder_5_io_a; // @[wallace.scala 54:25]
  wire  HalfAdder_5_io_b; // @[wallace.scala 54:25]
  wire  HalfAdder_5_io_s; // @[wallace.scala 54:25]
  wire  HalfAdder_5_io_co; // @[wallace.scala 54:25]
  wire  FullAdder_201_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_201_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_201_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_201_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_201_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_202_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_202_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_202_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_202_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_202_io_co; // @[wallace.scala 63:25]
  wire  FullAdder_203_io_a; // @[wallace.scala 63:25]
  wire  FullAdder_203_io_b; // @[wallace.scala 63:25]
  wire  FullAdder_203_io_ci; // @[wallace.scala 63:25]
  wire  FullAdder_203_io_s; // @[wallace.scala 63:25]
  wire  FullAdder_203_io_co; // @[wallace.scala 63:25]
  wire  res0_0 = io_pp_0[0]; // @[wallace.scala 34:43]
  wire  res0_1 = io_pp_0[1]; // @[wallace.scala 34:43]
  wire  res1_1 = io_pp_1[0]; // @[wallace.scala 34:43]
  wire  res0_30 = io_pp_15[15]; // @[wallace.scala 34:43]
  wire  res0_29 = FullAdder_75_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_28 = FullAdder_125_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_27 = FullAdder_157_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_26 = FullAdder_158_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_25 = FullAdder_179_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_24 = FullAdder_180_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_23 = FullAdder_181_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_22 = FullAdder_182_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_21 = FullAdder_195_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire [9:0] _T_264 = {res0_30,res0_29,res0_28,res0_27,res0_26,res0_25,res0_24,res0_23,res0_22,res0_21}; // @[Cat.scala 29:58]
  wire  res0_20 = FullAdder_196_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_19 = FullAdder_197_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_18 = FullAdder_198_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_17 = FullAdder_199_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_16 = FullAdder_200_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_15 = HalfAdder_3_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_14 = HalfAdder_4_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_13 = HalfAdder_5_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_12 = FullAdder_201_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire [18:0] _T_273 = {_T_264,res0_20,res0_19,res0_18,res0_17,res0_16,res0_15,res0_14,res0_13,res0_12}; // @[Cat.scala 29:58]
  wire  res0_11 = FullAdder_192_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_10 = FullAdder_202_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_9 = FullAdder_193_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_8 = FullAdder_177_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_7 = FullAdder_203_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_6 = FullAdder_194_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_5 = FullAdder_178_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_4 = FullAdder_156_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire  res0_3 = FullAdder_124_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire [27:0] _T_282 = {_T_273,res0_11,res0_10,res0_9,res0_8,res0_7,res0_6,res0_5,res0_4,res0_3}; // @[Cat.scala 29:58]
  wire  res0_2 = FullAdder_74_io_s; // @[wallace.scala 74:49 wallace.scala 79:13]
  wire [30:0] _T_285 = {_T_282,res0_2,res0_1,res0_0}; // @[Cat.scala 29:58]
  wire  res1_30 = FullAdder_75_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_29 = FullAdder_125_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_28 = FullAdder_157_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_27 = FullAdder_158_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_26 = FullAdder_179_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_25 = FullAdder_180_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_24 = FullAdder_181_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_23 = FullAdder_182_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_22 = FullAdder_195_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_21 = FullAdder_196_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire [9:0] _T_294 = {res1_30,res1_29,res1_28,res1_27,res1_26,res1_25,res1_24,res1_23,res1_22,res1_21}; // @[Cat.scala 29:58]
  wire  res1_20 = FullAdder_197_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_19 = FullAdder_198_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_18 = FullAdder_199_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_17 = FullAdder_200_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_16 = HalfAdder_3_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_15 = HalfAdder_4_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_14 = HalfAdder_5_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_13 = FullAdder_201_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire [18:0] _T_303 = {_T_294,res1_20,res1_19,res1_18,res1_17,res1_16,res1_15,res1_14,res1_13,1'h0}; // @[Cat.scala 29:58]
  wire  res1_11 = FullAdder_202_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire  res1_8 = FullAdder_203_io_co; // @[wallace.scala 75:49 wallace.scala 83:15]
  wire [27:0] _T_312 = {_T_303,res1_11,1'h0,1'h0,res1_8,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire [30:0] _T_315 = {_T_312,1'h0,res1_1,1'h0}; // @[Cat.scala 29:58]
  FullAdder FullAdder ( // @[wallace.scala 63:25]
    .io_a(FullAdder_io_a),
    .io_b(FullAdder_io_b),
    .io_ci(FullAdder_io_ci),
    .io_s(FullAdder_io_s),
    .io_co(FullAdder_io_co)
  );
  FullAdder FullAdder_1 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_1_io_a),
    .io_b(FullAdder_1_io_b),
    .io_ci(FullAdder_1_io_ci),
    .io_s(FullAdder_1_io_s),
    .io_co(FullAdder_1_io_co)
  );
  FullAdder FullAdder_2 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_2_io_a),
    .io_b(FullAdder_2_io_b),
    .io_ci(FullAdder_2_io_ci),
    .io_s(FullAdder_2_io_s),
    .io_co(FullAdder_2_io_co)
  );
  FullAdder FullAdder_3 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_3_io_a),
    .io_b(FullAdder_3_io_b),
    .io_ci(FullAdder_3_io_ci),
    .io_s(FullAdder_3_io_s),
    .io_co(FullAdder_3_io_co)
  );
  FullAdder FullAdder_4 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_4_io_a),
    .io_b(FullAdder_4_io_b),
    .io_ci(FullAdder_4_io_ci),
    .io_s(FullAdder_4_io_s),
    .io_co(FullAdder_4_io_co)
  );
  FullAdder FullAdder_5 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_5_io_a),
    .io_b(FullAdder_5_io_b),
    .io_ci(FullAdder_5_io_ci),
    .io_s(FullAdder_5_io_s),
    .io_co(FullAdder_5_io_co)
  );
  FullAdder FullAdder_6 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_6_io_a),
    .io_b(FullAdder_6_io_b),
    .io_ci(FullAdder_6_io_ci),
    .io_s(FullAdder_6_io_s),
    .io_co(FullAdder_6_io_co)
  );
  FullAdder FullAdder_7 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_7_io_a),
    .io_b(FullAdder_7_io_b),
    .io_ci(FullAdder_7_io_ci),
    .io_s(FullAdder_7_io_s),
    .io_co(FullAdder_7_io_co)
  );
  FullAdder FullAdder_8 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_8_io_a),
    .io_b(FullAdder_8_io_b),
    .io_ci(FullAdder_8_io_ci),
    .io_s(FullAdder_8_io_s),
    .io_co(FullAdder_8_io_co)
  );
  FullAdder FullAdder_9 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_9_io_a),
    .io_b(FullAdder_9_io_b),
    .io_ci(FullAdder_9_io_ci),
    .io_s(FullAdder_9_io_s),
    .io_co(FullAdder_9_io_co)
  );
  FullAdder FullAdder_10 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_10_io_a),
    .io_b(FullAdder_10_io_b),
    .io_ci(FullAdder_10_io_ci),
    .io_s(FullAdder_10_io_s),
    .io_co(FullAdder_10_io_co)
  );
  FullAdder FullAdder_11 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_11_io_a),
    .io_b(FullAdder_11_io_b),
    .io_ci(FullAdder_11_io_ci),
    .io_s(FullAdder_11_io_s),
    .io_co(FullAdder_11_io_co)
  );
  FullAdder FullAdder_12 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_12_io_a),
    .io_b(FullAdder_12_io_b),
    .io_ci(FullAdder_12_io_ci),
    .io_s(FullAdder_12_io_s),
    .io_co(FullAdder_12_io_co)
  );
  FullAdder FullAdder_13 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_13_io_a),
    .io_b(FullAdder_13_io_b),
    .io_ci(FullAdder_13_io_ci),
    .io_s(FullAdder_13_io_s),
    .io_co(FullAdder_13_io_co)
  );
  FullAdder FullAdder_14 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_14_io_a),
    .io_b(FullAdder_14_io_b),
    .io_ci(FullAdder_14_io_ci),
    .io_s(FullAdder_14_io_s),
    .io_co(FullAdder_14_io_co)
  );
  FullAdder FullAdder_15 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_15_io_a),
    .io_b(FullAdder_15_io_b),
    .io_ci(FullAdder_15_io_ci),
    .io_s(FullAdder_15_io_s),
    .io_co(FullAdder_15_io_co)
  );
  FullAdder FullAdder_16 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_16_io_a),
    .io_b(FullAdder_16_io_b),
    .io_ci(FullAdder_16_io_ci),
    .io_s(FullAdder_16_io_s),
    .io_co(FullAdder_16_io_co)
  );
  FullAdder FullAdder_17 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_17_io_a),
    .io_b(FullAdder_17_io_b),
    .io_ci(FullAdder_17_io_ci),
    .io_s(FullAdder_17_io_s),
    .io_co(FullAdder_17_io_co)
  );
  FullAdder FullAdder_18 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_18_io_a),
    .io_b(FullAdder_18_io_b),
    .io_ci(FullAdder_18_io_ci),
    .io_s(FullAdder_18_io_s),
    .io_co(FullAdder_18_io_co)
  );
  FullAdder FullAdder_19 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_19_io_a),
    .io_b(FullAdder_19_io_b),
    .io_ci(FullAdder_19_io_ci),
    .io_s(FullAdder_19_io_s),
    .io_co(FullAdder_19_io_co)
  );
  FullAdder FullAdder_20 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_20_io_a),
    .io_b(FullAdder_20_io_b),
    .io_ci(FullAdder_20_io_ci),
    .io_s(FullAdder_20_io_s),
    .io_co(FullAdder_20_io_co)
  );
  FullAdder FullAdder_21 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_21_io_a),
    .io_b(FullAdder_21_io_b),
    .io_ci(FullAdder_21_io_ci),
    .io_s(FullAdder_21_io_s),
    .io_co(FullAdder_21_io_co)
  );
  FullAdder FullAdder_22 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_22_io_a),
    .io_b(FullAdder_22_io_b),
    .io_ci(FullAdder_22_io_ci),
    .io_s(FullAdder_22_io_s),
    .io_co(FullAdder_22_io_co)
  );
  FullAdder FullAdder_23 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_23_io_a),
    .io_b(FullAdder_23_io_b),
    .io_ci(FullAdder_23_io_ci),
    .io_s(FullAdder_23_io_s),
    .io_co(FullAdder_23_io_co)
  );
  FullAdder FullAdder_24 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_24_io_a),
    .io_b(FullAdder_24_io_b),
    .io_ci(FullAdder_24_io_ci),
    .io_s(FullAdder_24_io_s),
    .io_co(FullAdder_24_io_co)
  );
  FullAdder FullAdder_25 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_25_io_a),
    .io_b(FullAdder_25_io_b),
    .io_ci(FullAdder_25_io_ci),
    .io_s(FullAdder_25_io_s),
    .io_co(FullAdder_25_io_co)
  );
  FullAdder FullAdder_26 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_26_io_a),
    .io_b(FullAdder_26_io_b),
    .io_ci(FullAdder_26_io_ci),
    .io_s(FullAdder_26_io_s),
    .io_co(FullAdder_26_io_co)
  );
  FullAdder FullAdder_27 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_27_io_a),
    .io_b(FullAdder_27_io_b),
    .io_ci(FullAdder_27_io_ci),
    .io_s(FullAdder_27_io_s),
    .io_co(FullAdder_27_io_co)
  );
  FullAdder FullAdder_28 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_28_io_a),
    .io_b(FullAdder_28_io_b),
    .io_ci(FullAdder_28_io_ci),
    .io_s(FullAdder_28_io_s),
    .io_co(FullAdder_28_io_co)
  );
  FullAdder FullAdder_29 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_29_io_a),
    .io_b(FullAdder_29_io_b),
    .io_ci(FullAdder_29_io_ci),
    .io_s(FullAdder_29_io_s),
    .io_co(FullAdder_29_io_co)
  );
  FullAdder FullAdder_30 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_30_io_a),
    .io_b(FullAdder_30_io_b),
    .io_ci(FullAdder_30_io_ci),
    .io_s(FullAdder_30_io_s),
    .io_co(FullAdder_30_io_co)
  );
  FullAdder FullAdder_31 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_31_io_a),
    .io_b(FullAdder_31_io_b),
    .io_ci(FullAdder_31_io_ci),
    .io_s(FullAdder_31_io_s),
    .io_co(FullAdder_31_io_co)
  );
  FullAdder FullAdder_32 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_32_io_a),
    .io_b(FullAdder_32_io_b),
    .io_ci(FullAdder_32_io_ci),
    .io_s(FullAdder_32_io_s),
    .io_co(FullAdder_32_io_co)
  );
  FullAdder FullAdder_33 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_33_io_a),
    .io_b(FullAdder_33_io_b),
    .io_ci(FullAdder_33_io_ci),
    .io_s(FullAdder_33_io_s),
    .io_co(FullAdder_33_io_co)
  );
  FullAdder FullAdder_34 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_34_io_a),
    .io_b(FullAdder_34_io_b),
    .io_ci(FullAdder_34_io_ci),
    .io_s(FullAdder_34_io_s),
    .io_co(FullAdder_34_io_co)
  );
  FullAdder FullAdder_35 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_35_io_a),
    .io_b(FullAdder_35_io_b),
    .io_ci(FullAdder_35_io_ci),
    .io_s(FullAdder_35_io_s),
    .io_co(FullAdder_35_io_co)
  );
  FullAdder FullAdder_36 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_36_io_a),
    .io_b(FullAdder_36_io_b),
    .io_ci(FullAdder_36_io_ci),
    .io_s(FullAdder_36_io_s),
    .io_co(FullAdder_36_io_co)
  );
  FullAdder FullAdder_37 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_37_io_a),
    .io_b(FullAdder_37_io_b),
    .io_ci(FullAdder_37_io_ci),
    .io_s(FullAdder_37_io_s),
    .io_co(FullAdder_37_io_co)
  );
  FullAdder FullAdder_38 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_38_io_a),
    .io_b(FullAdder_38_io_b),
    .io_ci(FullAdder_38_io_ci),
    .io_s(FullAdder_38_io_s),
    .io_co(FullAdder_38_io_co)
  );
  FullAdder FullAdder_39 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_39_io_a),
    .io_b(FullAdder_39_io_b),
    .io_ci(FullAdder_39_io_ci),
    .io_s(FullAdder_39_io_s),
    .io_co(FullAdder_39_io_co)
  );
  FullAdder FullAdder_40 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_40_io_a),
    .io_b(FullAdder_40_io_b),
    .io_ci(FullAdder_40_io_ci),
    .io_s(FullAdder_40_io_s),
    .io_co(FullAdder_40_io_co)
  );
  FullAdder FullAdder_41 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_41_io_a),
    .io_b(FullAdder_41_io_b),
    .io_ci(FullAdder_41_io_ci),
    .io_s(FullAdder_41_io_s),
    .io_co(FullAdder_41_io_co)
  );
  FullAdder FullAdder_42 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_42_io_a),
    .io_b(FullAdder_42_io_b),
    .io_ci(FullAdder_42_io_ci),
    .io_s(FullAdder_42_io_s),
    .io_co(FullAdder_42_io_co)
  );
  FullAdder FullAdder_43 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_43_io_a),
    .io_b(FullAdder_43_io_b),
    .io_ci(FullAdder_43_io_ci),
    .io_s(FullAdder_43_io_s),
    .io_co(FullAdder_43_io_co)
  );
  FullAdder FullAdder_44 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_44_io_a),
    .io_b(FullAdder_44_io_b),
    .io_ci(FullAdder_44_io_ci),
    .io_s(FullAdder_44_io_s),
    .io_co(FullAdder_44_io_co)
  );
  FullAdder FullAdder_45 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_45_io_a),
    .io_b(FullAdder_45_io_b),
    .io_ci(FullAdder_45_io_ci),
    .io_s(FullAdder_45_io_s),
    .io_co(FullAdder_45_io_co)
  );
  FullAdder FullAdder_46 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_46_io_a),
    .io_b(FullAdder_46_io_b),
    .io_ci(FullAdder_46_io_ci),
    .io_s(FullAdder_46_io_s),
    .io_co(FullAdder_46_io_co)
  );
  FullAdder FullAdder_47 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_47_io_a),
    .io_b(FullAdder_47_io_b),
    .io_ci(FullAdder_47_io_ci),
    .io_s(FullAdder_47_io_s),
    .io_co(FullAdder_47_io_co)
  );
  FullAdder FullAdder_48 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_48_io_a),
    .io_b(FullAdder_48_io_b),
    .io_ci(FullAdder_48_io_ci),
    .io_s(FullAdder_48_io_s),
    .io_co(FullAdder_48_io_co)
  );
  FullAdder FullAdder_49 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_49_io_a),
    .io_b(FullAdder_49_io_b),
    .io_ci(FullAdder_49_io_ci),
    .io_s(FullAdder_49_io_s),
    .io_co(FullAdder_49_io_co)
  );
  FullAdder FullAdder_50 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_50_io_a),
    .io_b(FullAdder_50_io_b),
    .io_ci(FullAdder_50_io_ci),
    .io_s(FullAdder_50_io_s),
    .io_co(FullAdder_50_io_co)
  );
  FullAdder FullAdder_51 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_51_io_a),
    .io_b(FullAdder_51_io_b),
    .io_ci(FullAdder_51_io_ci),
    .io_s(FullAdder_51_io_s),
    .io_co(FullAdder_51_io_co)
  );
  FullAdder FullAdder_52 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_52_io_a),
    .io_b(FullAdder_52_io_b),
    .io_ci(FullAdder_52_io_ci),
    .io_s(FullAdder_52_io_s),
    .io_co(FullAdder_52_io_co)
  );
  FullAdder FullAdder_53 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_53_io_a),
    .io_b(FullAdder_53_io_b),
    .io_ci(FullAdder_53_io_ci),
    .io_s(FullAdder_53_io_s),
    .io_co(FullAdder_53_io_co)
  );
  FullAdder FullAdder_54 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_54_io_a),
    .io_b(FullAdder_54_io_b),
    .io_ci(FullAdder_54_io_ci),
    .io_s(FullAdder_54_io_s),
    .io_co(FullAdder_54_io_co)
  );
  FullAdder FullAdder_55 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_55_io_a),
    .io_b(FullAdder_55_io_b),
    .io_ci(FullAdder_55_io_ci),
    .io_s(FullAdder_55_io_s),
    .io_co(FullAdder_55_io_co)
  );
  FullAdder FullAdder_56 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_56_io_a),
    .io_b(FullAdder_56_io_b),
    .io_ci(FullAdder_56_io_ci),
    .io_s(FullAdder_56_io_s),
    .io_co(FullAdder_56_io_co)
  );
  FullAdder FullAdder_57 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_57_io_a),
    .io_b(FullAdder_57_io_b),
    .io_ci(FullAdder_57_io_ci),
    .io_s(FullAdder_57_io_s),
    .io_co(FullAdder_57_io_co)
  );
  FullAdder FullAdder_58 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_58_io_a),
    .io_b(FullAdder_58_io_b),
    .io_ci(FullAdder_58_io_ci),
    .io_s(FullAdder_58_io_s),
    .io_co(FullAdder_58_io_co)
  );
  FullAdder FullAdder_59 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_59_io_a),
    .io_b(FullAdder_59_io_b),
    .io_ci(FullAdder_59_io_ci),
    .io_s(FullAdder_59_io_s),
    .io_co(FullAdder_59_io_co)
  );
  FullAdder FullAdder_60 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_60_io_a),
    .io_b(FullAdder_60_io_b),
    .io_ci(FullAdder_60_io_ci),
    .io_s(FullAdder_60_io_s),
    .io_co(FullAdder_60_io_co)
  );
  FullAdder FullAdder_61 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_61_io_a),
    .io_b(FullAdder_61_io_b),
    .io_ci(FullAdder_61_io_ci),
    .io_s(FullAdder_61_io_s),
    .io_co(FullAdder_61_io_co)
  );
  FullAdder FullAdder_62 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_62_io_a),
    .io_b(FullAdder_62_io_b),
    .io_ci(FullAdder_62_io_ci),
    .io_s(FullAdder_62_io_s),
    .io_co(FullAdder_62_io_co)
  );
  FullAdder FullAdder_63 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_63_io_a),
    .io_b(FullAdder_63_io_b),
    .io_ci(FullAdder_63_io_ci),
    .io_s(FullAdder_63_io_s),
    .io_co(FullAdder_63_io_co)
  );
  FullAdder FullAdder_64 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_64_io_a),
    .io_b(FullAdder_64_io_b),
    .io_ci(FullAdder_64_io_ci),
    .io_s(FullAdder_64_io_s),
    .io_co(FullAdder_64_io_co)
  );
  FullAdder FullAdder_65 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_65_io_a),
    .io_b(FullAdder_65_io_b),
    .io_ci(FullAdder_65_io_ci),
    .io_s(FullAdder_65_io_s),
    .io_co(FullAdder_65_io_co)
  );
  FullAdder FullAdder_66 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_66_io_a),
    .io_b(FullAdder_66_io_b),
    .io_ci(FullAdder_66_io_ci),
    .io_s(FullAdder_66_io_s),
    .io_co(FullAdder_66_io_co)
  );
  FullAdder FullAdder_67 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_67_io_a),
    .io_b(FullAdder_67_io_b),
    .io_ci(FullAdder_67_io_ci),
    .io_s(FullAdder_67_io_s),
    .io_co(FullAdder_67_io_co)
  );
  FullAdder FullAdder_68 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_68_io_a),
    .io_b(FullAdder_68_io_b),
    .io_ci(FullAdder_68_io_ci),
    .io_s(FullAdder_68_io_s),
    .io_co(FullAdder_68_io_co)
  );
  FullAdder FullAdder_69 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_69_io_a),
    .io_b(FullAdder_69_io_b),
    .io_ci(FullAdder_69_io_ci),
    .io_s(FullAdder_69_io_s),
    .io_co(FullAdder_69_io_co)
  );
  FullAdder FullAdder_70 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_70_io_a),
    .io_b(FullAdder_70_io_b),
    .io_ci(FullAdder_70_io_ci),
    .io_s(FullAdder_70_io_s),
    .io_co(FullAdder_70_io_co)
  );
  FullAdder FullAdder_71 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_71_io_a),
    .io_b(FullAdder_71_io_b),
    .io_ci(FullAdder_71_io_ci),
    .io_s(FullAdder_71_io_s),
    .io_co(FullAdder_71_io_co)
  );
  FullAdder FullAdder_72 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_72_io_a),
    .io_b(FullAdder_72_io_b),
    .io_ci(FullAdder_72_io_ci),
    .io_s(FullAdder_72_io_s),
    .io_co(FullAdder_72_io_co)
  );
  FullAdder FullAdder_73 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_73_io_a),
    .io_b(FullAdder_73_io_b),
    .io_ci(FullAdder_73_io_ci),
    .io_s(FullAdder_73_io_s),
    .io_co(FullAdder_73_io_co)
  );
  FullAdder FullAdder_74 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_74_io_a),
    .io_b(FullAdder_74_io_b),
    .io_ci(FullAdder_74_io_ci),
    .io_s(FullAdder_74_io_s),
    .io_co(FullAdder_74_io_co)
  );
  FullAdder FullAdder_75 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_75_io_a),
    .io_b(FullAdder_75_io_b),
    .io_ci(FullAdder_75_io_ci),
    .io_s(FullAdder_75_io_s),
    .io_co(FullAdder_75_io_co)
  );
  FullAdder FullAdder_76 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_76_io_a),
    .io_b(FullAdder_76_io_b),
    .io_ci(FullAdder_76_io_ci),
    .io_s(FullAdder_76_io_s),
    .io_co(FullAdder_76_io_co)
  );
  FullAdder FullAdder_77 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_77_io_a),
    .io_b(FullAdder_77_io_b),
    .io_ci(FullAdder_77_io_ci),
    .io_s(FullAdder_77_io_s),
    .io_co(FullAdder_77_io_co)
  );
  FullAdder FullAdder_78 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_78_io_a),
    .io_b(FullAdder_78_io_b),
    .io_ci(FullAdder_78_io_ci),
    .io_s(FullAdder_78_io_s),
    .io_co(FullAdder_78_io_co)
  );
  FullAdder FullAdder_79 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_79_io_a),
    .io_b(FullAdder_79_io_b),
    .io_ci(FullAdder_79_io_ci),
    .io_s(FullAdder_79_io_s),
    .io_co(FullAdder_79_io_co)
  );
  FullAdder FullAdder_80 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_80_io_a),
    .io_b(FullAdder_80_io_b),
    .io_ci(FullAdder_80_io_ci),
    .io_s(FullAdder_80_io_s),
    .io_co(FullAdder_80_io_co)
  );
  FullAdder FullAdder_81 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_81_io_a),
    .io_b(FullAdder_81_io_b),
    .io_ci(FullAdder_81_io_ci),
    .io_s(FullAdder_81_io_s),
    .io_co(FullAdder_81_io_co)
  );
  FullAdder FullAdder_82 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_82_io_a),
    .io_b(FullAdder_82_io_b),
    .io_ci(FullAdder_82_io_ci),
    .io_s(FullAdder_82_io_s),
    .io_co(FullAdder_82_io_co)
  );
  FullAdder FullAdder_83 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_83_io_a),
    .io_b(FullAdder_83_io_b),
    .io_ci(FullAdder_83_io_ci),
    .io_s(FullAdder_83_io_s),
    .io_co(FullAdder_83_io_co)
  );
  FullAdder FullAdder_84 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_84_io_a),
    .io_b(FullAdder_84_io_b),
    .io_ci(FullAdder_84_io_ci),
    .io_s(FullAdder_84_io_s),
    .io_co(FullAdder_84_io_co)
  );
  FullAdder FullAdder_85 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_85_io_a),
    .io_b(FullAdder_85_io_b),
    .io_ci(FullAdder_85_io_ci),
    .io_s(FullAdder_85_io_s),
    .io_co(FullAdder_85_io_co)
  );
  FullAdder FullAdder_86 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_86_io_a),
    .io_b(FullAdder_86_io_b),
    .io_ci(FullAdder_86_io_ci),
    .io_s(FullAdder_86_io_s),
    .io_co(FullAdder_86_io_co)
  );
  FullAdder FullAdder_87 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_87_io_a),
    .io_b(FullAdder_87_io_b),
    .io_ci(FullAdder_87_io_ci),
    .io_s(FullAdder_87_io_s),
    .io_co(FullAdder_87_io_co)
  );
  FullAdder FullAdder_88 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_88_io_a),
    .io_b(FullAdder_88_io_b),
    .io_ci(FullAdder_88_io_ci),
    .io_s(FullAdder_88_io_s),
    .io_co(FullAdder_88_io_co)
  );
  FullAdder FullAdder_89 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_89_io_a),
    .io_b(FullAdder_89_io_b),
    .io_ci(FullAdder_89_io_ci),
    .io_s(FullAdder_89_io_s),
    .io_co(FullAdder_89_io_co)
  );
  FullAdder FullAdder_90 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_90_io_a),
    .io_b(FullAdder_90_io_b),
    .io_ci(FullAdder_90_io_ci),
    .io_s(FullAdder_90_io_s),
    .io_co(FullAdder_90_io_co)
  );
  FullAdder FullAdder_91 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_91_io_a),
    .io_b(FullAdder_91_io_b),
    .io_ci(FullAdder_91_io_ci),
    .io_s(FullAdder_91_io_s),
    .io_co(FullAdder_91_io_co)
  );
  FullAdder FullAdder_92 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_92_io_a),
    .io_b(FullAdder_92_io_b),
    .io_ci(FullAdder_92_io_ci),
    .io_s(FullAdder_92_io_s),
    .io_co(FullAdder_92_io_co)
  );
  FullAdder FullAdder_93 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_93_io_a),
    .io_b(FullAdder_93_io_b),
    .io_ci(FullAdder_93_io_ci),
    .io_s(FullAdder_93_io_s),
    .io_co(FullAdder_93_io_co)
  );
  FullAdder FullAdder_94 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_94_io_a),
    .io_b(FullAdder_94_io_b),
    .io_ci(FullAdder_94_io_ci),
    .io_s(FullAdder_94_io_s),
    .io_co(FullAdder_94_io_co)
  );
  FullAdder FullAdder_95 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_95_io_a),
    .io_b(FullAdder_95_io_b),
    .io_ci(FullAdder_95_io_ci),
    .io_s(FullAdder_95_io_s),
    .io_co(FullAdder_95_io_co)
  );
  FullAdder FullAdder_96 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_96_io_a),
    .io_b(FullAdder_96_io_b),
    .io_ci(FullAdder_96_io_ci),
    .io_s(FullAdder_96_io_s),
    .io_co(FullAdder_96_io_co)
  );
  FullAdder FullAdder_97 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_97_io_a),
    .io_b(FullAdder_97_io_b),
    .io_ci(FullAdder_97_io_ci),
    .io_s(FullAdder_97_io_s),
    .io_co(FullAdder_97_io_co)
  );
  FullAdder FullAdder_98 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_98_io_a),
    .io_b(FullAdder_98_io_b),
    .io_ci(FullAdder_98_io_ci),
    .io_s(FullAdder_98_io_s),
    .io_co(FullAdder_98_io_co)
  );
  FullAdder FullAdder_99 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_99_io_a),
    .io_b(FullAdder_99_io_b),
    .io_ci(FullAdder_99_io_ci),
    .io_s(FullAdder_99_io_s),
    .io_co(FullAdder_99_io_co)
  );
  FullAdder FullAdder_100 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_100_io_a),
    .io_b(FullAdder_100_io_b),
    .io_ci(FullAdder_100_io_ci),
    .io_s(FullAdder_100_io_s),
    .io_co(FullAdder_100_io_co)
  );
  FullAdder FullAdder_101 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_101_io_a),
    .io_b(FullAdder_101_io_b),
    .io_ci(FullAdder_101_io_ci),
    .io_s(FullAdder_101_io_s),
    .io_co(FullAdder_101_io_co)
  );
  FullAdder FullAdder_102 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_102_io_a),
    .io_b(FullAdder_102_io_b),
    .io_ci(FullAdder_102_io_ci),
    .io_s(FullAdder_102_io_s),
    .io_co(FullAdder_102_io_co)
  );
  FullAdder FullAdder_103 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_103_io_a),
    .io_b(FullAdder_103_io_b),
    .io_ci(FullAdder_103_io_ci),
    .io_s(FullAdder_103_io_s),
    .io_co(FullAdder_103_io_co)
  );
  FullAdder FullAdder_104 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_104_io_a),
    .io_b(FullAdder_104_io_b),
    .io_ci(FullAdder_104_io_ci),
    .io_s(FullAdder_104_io_s),
    .io_co(FullAdder_104_io_co)
  );
  FullAdder FullAdder_105 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_105_io_a),
    .io_b(FullAdder_105_io_b),
    .io_ci(FullAdder_105_io_ci),
    .io_s(FullAdder_105_io_s),
    .io_co(FullAdder_105_io_co)
  );
  FullAdder FullAdder_106 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_106_io_a),
    .io_b(FullAdder_106_io_b),
    .io_ci(FullAdder_106_io_ci),
    .io_s(FullAdder_106_io_s),
    .io_co(FullAdder_106_io_co)
  );
  FullAdder FullAdder_107 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_107_io_a),
    .io_b(FullAdder_107_io_b),
    .io_ci(FullAdder_107_io_ci),
    .io_s(FullAdder_107_io_s),
    .io_co(FullAdder_107_io_co)
  );
  FullAdder FullAdder_108 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_108_io_a),
    .io_b(FullAdder_108_io_b),
    .io_ci(FullAdder_108_io_ci),
    .io_s(FullAdder_108_io_s),
    .io_co(FullAdder_108_io_co)
  );
  FullAdder FullAdder_109 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_109_io_a),
    .io_b(FullAdder_109_io_b),
    .io_ci(FullAdder_109_io_ci),
    .io_s(FullAdder_109_io_s),
    .io_co(FullAdder_109_io_co)
  );
  FullAdder FullAdder_110 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_110_io_a),
    .io_b(FullAdder_110_io_b),
    .io_ci(FullAdder_110_io_ci),
    .io_s(FullAdder_110_io_s),
    .io_co(FullAdder_110_io_co)
  );
  FullAdder FullAdder_111 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_111_io_a),
    .io_b(FullAdder_111_io_b),
    .io_ci(FullAdder_111_io_ci),
    .io_s(FullAdder_111_io_s),
    .io_co(FullAdder_111_io_co)
  );
  FullAdder FullAdder_112 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_112_io_a),
    .io_b(FullAdder_112_io_b),
    .io_ci(FullAdder_112_io_ci),
    .io_s(FullAdder_112_io_s),
    .io_co(FullAdder_112_io_co)
  );
  FullAdder FullAdder_113 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_113_io_a),
    .io_b(FullAdder_113_io_b),
    .io_ci(FullAdder_113_io_ci),
    .io_s(FullAdder_113_io_s),
    .io_co(FullAdder_113_io_co)
  );
  FullAdder FullAdder_114 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_114_io_a),
    .io_b(FullAdder_114_io_b),
    .io_ci(FullAdder_114_io_ci),
    .io_s(FullAdder_114_io_s),
    .io_co(FullAdder_114_io_co)
  );
  FullAdder FullAdder_115 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_115_io_a),
    .io_b(FullAdder_115_io_b),
    .io_ci(FullAdder_115_io_ci),
    .io_s(FullAdder_115_io_s),
    .io_co(FullAdder_115_io_co)
  );
  FullAdder FullAdder_116 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_116_io_a),
    .io_b(FullAdder_116_io_b),
    .io_ci(FullAdder_116_io_ci),
    .io_s(FullAdder_116_io_s),
    .io_co(FullAdder_116_io_co)
  );
  FullAdder FullAdder_117 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_117_io_a),
    .io_b(FullAdder_117_io_b),
    .io_ci(FullAdder_117_io_ci),
    .io_s(FullAdder_117_io_s),
    .io_co(FullAdder_117_io_co)
  );
  FullAdder FullAdder_118 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_118_io_a),
    .io_b(FullAdder_118_io_b),
    .io_ci(FullAdder_118_io_ci),
    .io_s(FullAdder_118_io_s),
    .io_co(FullAdder_118_io_co)
  );
  FullAdder FullAdder_119 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_119_io_a),
    .io_b(FullAdder_119_io_b),
    .io_ci(FullAdder_119_io_ci),
    .io_s(FullAdder_119_io_s),
    .io_co(FullAdder_119_io_co)
  );
  FullAdder FullAdder_120 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_120_io_a),
    .io_b(FullAdder_120_io_b),
    .io_ci(FullAdder_120_io_ci),
    .io_s(FullAdder_120_io_s),
    .io_co(FullAdder_120_io_co)
  );
  FullAdder FullAdder_121 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_121_io_a),
    .io_b(FullAdder_121_io_b),
    .io_ci(FullAdder_121_io_ci),
    .io_s(FullAdder_121_io_s),
    .io_co(FullAdder_121_io_co)
  );
  FullAdder FullAdder_122 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_122_io_a),
    .io_b(FullAdder_122_io_b),
    .io_ci(FullAdder_122_io_ci),
    .io_s(FullAdder_122_io_s),
    .io_co(FullAdder_122_io_co)
  );
  FullAdder FullAdder_123 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_123_io_a),
    .io_b(FullAdder_123_io_b),
    .io_ci(FullAdder_123_io_ci),
    .io_s(FullAdder_123_io_s),
    .io_co(FullAdder_123_io_co)
  );
  FullAdder FullAdder_124 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_124_io_a),
    .io_b(FullAdder_124_io_b),
    .io_ci(FullAdder_124_io_ci),
    .io_s(FullAdder_124_io_s),
    .io_co(FullAdder_124_io_co)
  );
  FullAdder FullAdder_125 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_125_io_a),
    .io_b(FullAdder_125_io_b),
    .io_ci(FullAdder_125_io_ci),
    .io_s(FullAdder_125_io_s),
    .io_co(FullAdder_125_io_co)
  );
  FullAdder FullAdder_126 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_126_io_a),
    .io_b(FullAdder_126_io_b),
    .io_ci(FullAdder_126_io_ci),
    .io_s(FullAdder_126_io_s),
    .io_co(FullAdder_126_io_co)
  );
  FullAdder FullAdder_127 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_127_io_a),
    .io_b(FullAdder_127_io_b),
    .io_ci(FullAdder_127_io_ci),
    .io_s(FullAdder_127_io_s),
    .io_co(FullAdder_127_io_co)
  );
  FullAdder FullAdder_128 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_128_io_a),
    .io_b(FullAdder_128_io_b),
    .io_ci(FullAdder_128_io_ci),
    .io_s(FullAdder_128_io_s),
    .io_co(FullAdder_128_io_co)
  );
  FullAdder FullAdder_129 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_129_io_a),
    .io_b(FullAdder_129_io_b),
    .io_ci(FullAdder_129_io_ci),
    .io_s(FullAdder_129_io_s),
    .io_co(FullAdder_129_io_co)
  );
  FullAdder FullAdder_130 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_130_io_a),
    .io_b(FullAdder_130_io_b),
    .io_ci(FullAdder_130_io_ci),
    .io_s(FullAdder_130_io_s),
    .io_co(FullAdder_130_io_co)
  );
  FullAdder FullAdder_131 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_131_io_a),
    .io_b(FullAdder_131_io_b),
    .io_ci(FullAdder_131_io_ci),
    .io_s(FullAdder_131_io_s),
    .io_co(FullAdder_131_io_co)
  );
  FullAdder FullAdder_132 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_132_io_a),
    .io_b(FullAdder_132_io_b),
    .io_ci(FullAdder_132_io_ci),
    .io_s(FullAdder_132_io_s),
    .io_co(FullAdder_132_io_co)
  );
  FullAdder FullAdder_133 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_133_io_a),
    .io_b(FullAdder_133_io_b),
    .io_ci(FullAdder_133_io_ci),
    .io_s(FullAdder_133_io_s),
    .io_co(FullAdder_133_io_co)
  );
  FullAdder FullAdder_134 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_134_io_a),
    .io_b(FullAdder_134_io_b),
    .io_ci(FullAdder_134_io_ci),
    .io_s(FullAdder_134_io_s),
    .io_co(FullAdder_134_io_co)
  );
  FullAdder FullAdder_135 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_135_io_a),
    .io_b(FullAdder_135_io_b),
    .io_ci(FullAdder_135_io_ci),
    .io_s(FullAdder_135_io_s),
    .io_co(FullAdder_135_io_co)
  );
  FullAdder FullAdder_136 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_136_io_a),
    .io_b(FullAdder_136_io_b),
    .io_ci(FullAdder_136_io_ci),
    .io_s(FullAdder_136_io_s),
    .io_co(FullAdder_136_io_co)
  );
  FullAdder FullAdder_137 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_137_io_a),
    .io_b(FullAdder_137_io_b),
    .io_ci(FullAdder_137_io_ci),
    .io_s(FullAdder_137_io_s),
    .io_co(FullAdder_137_io_co)
  );
  FullAdder FullAdder_138 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_138_io_a),
    .io_b(FullAdder_138_io_b),
    .io_ci(FullAdder_138_io_ci),
    .io_s(FullAdder_138_io_s),
    .io_co(FullAdder_138_io_co)
  );
  FullAdder FullAdder_139 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_139_io_a),
    .io_b(FullAdder_139_io_b),
    .io_ci(FullAdder_139_io_ci),
    .io_s(FullAdder_139_io_s),
    .io_co(FullAdder_139_io_co)
  );
  FullAdder FullAdder_140 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_140_io_a),
    .io_b(FullAdder_140_io_b),
    .io_ci(FullAdder_140_io_ci),
    .io_s(FullAdder_140_io_s),
    .io_co(FullAdder_140_io_co)
  );
  FullAdder FullAdder_141 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_141_io_a),
    .io_b(FullAdder_141_io_b),
    .io_ci(FullAdder_141_io_ci),
    .io_s(FullAdder_141_io_s),
    .io_co(FullAdder_141_io_co)
  );
  FullAdder FullAdder_142 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_142_io_a),
    .io_b(FullAdder_142_io_b),
    .io_ci(FullAdder_142_io_ci),
    .io_s(FullAdder_142_io_s),
    .io_co(FullAdder_142_io_co)
  );
  FullAdder FullAdder_143 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_143_io_a),
    .io_b(FullAdder_143_io_b),
    .io_ci(FullAdder_143_io_ci),
    .io_s(FullAdder_143_io_s),
    .io_co(FullAdder_143_io_co)
  );
  FullAdder FullAdder_144 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_144_io_a),
    .io_b(FullAdder_144_io_b),
    .io_ci(FullAdder_144_io_ci),
    .io_s(FullAdder_144_io_s),
    .io_co(FullAdder_144_io_co)
  );
  FullAdder FullAdder_145 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_145_io_a),
    .io_b(FullAdder_145_io_b),
    .io_ci(FullAdder_145_io_ci),
    .io_s(FullAdder_145_io_s),
    .io_co(FullAdder_145_io_co)
  );
  FullAdder FullAdder_146 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_146_io_a),
    .io_b(FullAdder_146_io_b),
    .io_ci(FullAdder_146_io_ci),
    .io_s(FullAdder_146_io_s),
    .io_co(FullAdder_146_io_co)
  );
  FullAdder FullAdder_147 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_147_io_a),
    .io_b(FullAdder_147_io_b),
    .io_ci(FullAdder_147_io_ci),
    .io_s(FullAdder_147_io_s),
    .io_co(FullAdder_147_io_co)
  );
  FullAdder FullAdder_148 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_148_io_a),
    .io_b(FullAdder_148_io_b),
    .io_ci(FullAdder_148_io_ci),
    .io_s(FullAdder_148_io_s),
    .io_co(FullAdder_148_io_co)
  );
  FullAdder FullAdder_149 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_149_io_a),
    .io_b(FullAdder_149_io_b),
    .io_ci(FullAdder_149_io_ci),
    .io_s(FullAdder_149_io_s),
    .io_co(FullAdder_149_io_co)
  );
  FullAdder FullAdder_150 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_150_io_a),
    .io_b(FullAdder_150_io_b),
    .io_ci(FullAdder_150_io_ci),
    .io_s(FullAdder_150_io_s),
    .io_co(FullAdder_150_io_co)
  );
  FullAdder FullAdder_151 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_151_io_a),
    .io_b(FullAdder_151_io_b),
    .io_ci(FullAdder_151_io_ci),
    .io_s(FullAdder_151_io_s),
    .io_co(FullAdder_151_io_co)
  );
  FullAdder FullAdder_152 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_152_io_a),
    .io_b(FullAdder_152_io_b),
    .io_ci(FullAdder_152_io_ci),
    .io_s(FullAdder_152_io_s),
    .io_co(FullAdder_152_io_co)
  );
  FullAdder FullAdder_153 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_153_io_a),
    .io_b(FullAdder_153_io_b),
    .io_ci(FullAdder_153_io_ci),
    .io_s(FullAdder_153_io_s),
    .io_co(FullAdder_153_io_co)
  );
  HalfAdder HalfAdder ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_io_a),
    .io_b(HalfAdder_io_b),
    .io_s(HalfAdder_io_s),
    .io_co(HalfAdder_io_co)
  );
  FullAdder FullAdder_154 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_154_io_a),
    .io_b(FullAdder_154_io_b),
    .io_ci(FullAdder_154_io_ci),
    .io_s(FullAdder_154_io_s),
    .io_co(FullAdder_154_io_co)
  );
  FullAdder FullAdder_155 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_155_io_a),
    .io_b(FullAdder_155_io_b),
    .io_ci(FullAdder_155_io_ci),
    .io_s(FullAdder_155_io_s),
    .io_co(FullAdder_155_io_co)
  );
  FullAdder FullAdder_156 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_156_io_a),
    .io_b(FullAdder_156_io_b),
    .io_ci(FullAdder_156_io_ci),
    .io_s(FullAdder_156_io_s),
    .io_co(FullAdder_156_io_co)
  );
  FullAdder FullAdder_157 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_157_io_a),
    .io_b(FullAdder_157_io_b),
    .io_ci(FullAdder_157_io_ci),
    .io_s(FullAdder_157_io_s),
    .io_co(FullAdder_157_io_co)
  );
  FullAdder FullAdder_158 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_158_io_a),
    .io_b(FullAdder_158_io_b),
    .io_ci(FullAdder_158_io_ci),
    .io_s(FullAdder_158_io_s),
    .io_co(FullAdder_158_io_co)
  );
  FullAdder FullAdder_159 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_159_io_a),
    .io_b(FullAdder_159_io_b),
    .io_ci(FullAdder_159_io_ci),
    .io_s(FullAdder_159_io_s),
    .io_co(FullAdder_159_io_co)
  );
  FullAdder FullAdder_160 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_160_io_a),
    .io_b(FullAdder_160_io_b),
    .io_ci(FullAdder_160_io_ci),
    .io_s(FullAdder_160_io_s),
    .io_co(FullAdder_160_io_co)
  );
  FullAdder FullAdder_161 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_161_io_a),
    .io_b(FullAdder_161_io_b),
    .io_ci(FullAdder_161_io_ci),
    .io_s(FullAdder_161_io_s),
    .io_co(FullAdder_161_io_co)
  );
  FullAdder FullAdder_162 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_162_io_a),
    .io_b(FullAdder_162_io_b),
    .io_ci(FullAdder_162_io_ci),
    .io_s(FullAdder_162_io_s),
    .io_co(FullAdder_162_io_co)
  );
  FullAdder FullAdder_163 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_163_io_a),
    .io_b(FullAdder_163_io_b),
    .io_ci(FullAdder_163_io_ci),
    .io_s(FullAdder_163_io_s),
    .io_co(FullAdder_163_io_co)
  );
  FullAdder FullAdder_164 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_164_io_a),
    .io_b(FullAdder_164_io_b),
    .io_ci(FullAdder_164_io_ci),
    .io_s(FullAdder_164_io_s),
    .io_co(FullAdder_164_io_co)
  );
  FullAdder FullAdder_165 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_165_io_a),
    .io_b(FullAdder_165_io_b),
    .io_ci(FullAdder_165_io_ci),
    .io_s(FullAdder_165_io_s),
    .io_co(FullAdder_165_io_co)
  );
  FullAdder FullAdder_166 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_166_io_a),
    .io_b(FullAdder_166_io_b),
    .io_ci(FullAdder_166_io_ci),
    .io_s(FullAdder_166_io_s),
    .io_co(FullAdder_166_io_co)
  );
  FullAdder FullAdder_167 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_167_io_a),
    .io_b(FullAdder_167_io_b),
    .io_ci(FullAdder_167_io_ci),
    .io_s(FullAdder_167_io_s),
    .io_co(FullAdder_167_io_co)
  );
  FullAdder FullAdder_168 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_168_io_a),
    .io_b(FullAdder_168_io_b),
    .io_ci(FullAdder_168_io_ci),
    .io_s(FullAdder_168_io_s),
    .io_co(FullAdder_168_io_co)
  );
  FullAdder FullAdder_169 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_169_io_a),
    .io_b(FullAdder_169_io_b),
    .io_ci(FullAdder_169_io_ci),
    .io_s(FullAdder_169_io_s),
    .io_co(FullAdder_169_io_co)
  );
  FullAdder FullAdder_170 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_170_io_a),
    .io_b(FullAdder_170_io_b),
    .io_ci(FullAdder_170_io_ci),
    .io_s(FullAdder_170_io_s),
    .io_co(FullAdder_170_io_co)
  );
  FullAdder FullAdder_171 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_171_io_a),
    .io_b(FullAdder_171_io_b),
    .io_ci(FullAdder_171_io_ci),
    .io_s(FullAdder_171_io_s),
    .io_co(FullAdder_171_io_co)
  );
  FullAdder FullAdder_172 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_172_io_a),
    .io_b(FullAdder_172_io_b),
    .io_ci(FullAdder_172_io_ci),
    .io_s(FullAdder_172_io_s),
    .io_co(FullAdder_172_io_co)
  );
  FullAdder FullAdder_173 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_173_io_a),
    .io_b(FullAdder_173_io_b),
    .io_ci(FullAdder_173_io_ci),
    .io_s(FullAdder_173_io_s),
    .io_co(FullAdder_173_io_co)
  );
  FullAdder FullAdder_174 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_174_io_a),
    .io_b(FullAdder_174_io_b),
    .io_ci(FullAdder_174_io_ci),
    .io_s(FullAdder_174_io_s),
    .io_co(FullAdder_174_io_co)
  );
  HalfAdder HalfAdder_1 ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_1_io_a),
    .io_b(HalfAdder_1_io_b),
    .io_s(HalfAdder_1_io_s),
    .io_co(HalfAdder_1_io_co)
  );
  FullAdder FullAdder_175 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_175_io_a),
    .io_b(FullAdder_175_io_b),
    .io_ci(FullAdder_175_io_ci),
    .io_s(FullAdder_175_io_s),
    .io_co(FullAdder_175_io_co)
  );
  FullAdder FullAdder_176 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_176_io_a),
    .io_b(FullAdder_176_io_b),
    .io_ci(FullAdder_176_io_ci),
    .io_s(FullAdder_176_io_s),
    .io_co(FullAdder_176_io_co)
  );
  FullAdder FullAdder_177 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_177_io_a),
    .io_b(FullAdder_177_io_b),
    .io_ci(FullAdder_177_io_ci),
    .io_s(FullAdder_177_io_s),
    .io_co(FullAdder_177_io_co)
  );
  FullAdder FullAdder_178 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_178_io_a),
    .io_b(FullAdder_178_io_b),
    .io_ci(FullAdder_178_io_ci),
    .io_s(FullAdder_178_io_s),
    .io_co(FullAdder_178_io_co)
  );
  FullAdder FullAdder_179 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_179_io_a),
    .io_b(FullAdder_179_io_b),
    .io_ci(FullAdder_179_io_ci),
    .io_s(FullAdder_179_io_s),
    .io_co(FullAdder_179_io_co)
  );
  FullAdder FullAdder_180 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_180_io_a),
    .io_b(FullAdder_180_io_b),
    .io_ci(FullAdder_180_io_ci),
    .io_s(FullAdder_180_io_s),
    .io_co(FullAdder_180_io_co)
  );
  FullAdder FullAdder_181 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_181_io_a),
    .io_b(FullAdder_181_io_b),
    .io_ci(FullAdder_181_io_ci),
    .io_s(FullAdder_181_io_s),
    .io_co(FullAdder_181_io_co)
  );
  FullAdder FullAdder_182 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_182_io_a),
    .io_b(FullAdder_182_io_b),
    .io_ci(FullAdder_182_io_ci),
    .io_s(FullAdder_182_io_s),
    .io_co(FullAdder_182_io_co)
  );
  FullAdder FullAdder_183 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_183_io_a),
    .io_b(FullAdder_183_io_b),
    .io_ci(FullAdder_183_io_ci),
    .io_s(FullAdder_183_io_s),
    .io_co(FullAdder_183_io_co)
  );
  FullAdder FullAdder_184 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_184_io_a),
    .io_b(FullAdder_184_io_b),
    .io_ci(FullAdder_184_io_ci),
    .io_s(FullAdder_184_io_s),
    .io_co(FullAdder_184_io_co)
  );
  FullAdder FullAdder_185 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_185_io_a),
    .io_b(FullAdder_185_io_b),
    .io_ci(FullAdder_185_io_ci),
    .io_s(FullAdder_185_io_s),
    .io_co(FullAdder_185_io_co)
  );
  FullAdder FullAdder_186 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_186_io_a),
    .io_b(FullAdder_186_io_b),
    .io_ci(FullAdder_186_io_ci),
    .io_s(FullAdder_186_io_s),
    .io_co(FullAdder_186_io_co)
  );
  FullAdder FullAdder_187 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_187_io_a),
    .io_b(FullAdder_187_io_b),
    .io_ci(FullAdder_187_io_ci),
    .io_s(FullAdder_187_io_s),
    .io_co(FullAdder_187_io_co)
  );
  HalfAdder HalfAdder_2 ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_2_io_a),
    .io_b(HalfAdder_2_io_b),
    .io_s(HalfAdder_2_io_s),
    .io_co(HalfAdder_2_io_co)
  );
  FullAdder FullAdder_188 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_188_io_a),
    .io_b(FullAdder_188_io_b),
    .io_ci(FullAdder_188_io_ci),
    .io_s(FullAdder_188_io_s),
    .io_co(FullAdder_188_io_co)
  );
  FullAdder FullAdder_189 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_189_io_a),
    .io_b(FullAdder_189_io_b),
    .io_ci(FullAdder_189_io_ci),
    .io_s(FullAdder_189_io_s),
    .io_co(FullAdder_189_io_co)
  );
  FullAdder FullAdder_190 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_190_io_a),
    .io_b(FullAdder_190_io_b),
    .io_ci(FullAdder_190_io_ci),
    .io_s(FullAdder_190_io_s),
    .io_co(FullAdder_190_io_co)
  );
  FullAdder FullAdder_191 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_191_io_a),
    .io_b(FullAdder_191_io_b),
    .io_ci(FullAdder_191_io_ci),
    .io_s(FullAdder_191_io_s),
    .io_co(FullAdder_191_io_co)
  );
  FullAdder FullAdder_192 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_192_io_a),
    .io_b(FullAdder_192_io_b),
    .io_ci(FullAdder_192_io_ci),
    .io_s(FullAdder_192_io_s),
    .io_co(FullAdder_192_io_co)
  );
  FullAdder FullAdder_193 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_193_io_a),
    .io_b(FullAdder_193_io_b),
    .io_ci(FullAdder_193_io_ci),
    .io_s(FullAdder_193_io_s),
    .io_co(FullAdder_193_io_co)
  );
  FullAdder FullAdder_194 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_194_io_a),
    .io_b(FullAdder_194_io_b),
    .io_ci(FullAdder_194_io_ci),
    .io_s(FullAdder_194_io_s),
    .io_co(FullAdder_194_io_co)
  );
  FullAdder FullAdder_195 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_195_io_a),
    .io_b(FullAdder_195_io_b),
    .io_ci(FullAdder_195_io_ci),
    .io_s(FullAdder_195_io_s),
    .io_co(FullAdder_195_io_co)
  );
  FullAdder FullAdder_196 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_196_io_a),
    .io_b(FullAdder_196_io_b),
    .io_ci(FullAdder_196_io_ci),
    .io_s(FullAdder_196_io_s),
    .io_co(FullAdder_196_io_co)
  );
  FullAdder FullAdder_197 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_197_io_a),
    .io_b(FullAdder_197_io_b),
    .io_ci(FullAdder_197_io_ci),
    .io_s(FullAdder_197_io_s),
    .io_co(FullAdder_197_io_co)
  );
  FullAdder FullAdder_198 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_198_io_a),
    .io_b(FullAdder_198_io_b),
    .io_ci(FullAdder_198_io_ci),
    .io_s(FullAdder_198_io_s),
    .io_co(FullAdder_198_io_co)
  );
  FullAdder FullAdder_199 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_199_io_a),
    .io_b(FullAdder_199_io_b),
    .io_ci(FullAdder_199_io_ci),
    .io_s(FullAdder_199_io_s),
    .io_co(FullAdder_199_io_co)
  );
  FullAdder FullAdder_200 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_200_io_a),
    .io_b(FullAdder_200_io_b),
    .io_ci(FullAdder_200_io_ci),
    .io_s(FullAdder_200_io_s),
    .io_co(FullAdder_200_io_co)
  );
  HalfAdder HalfAdder_3 ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_3_io_a),
    .io_b(HalfAdder_3_io_b),
    .io_s(HalfAdder_3_io_s),
    .io_co(HalfAdder_3_io_co)
  );
  HalfAdder HalfAdder_4 ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_4_io_a),
    .io_b(HalfAdder_4_io_b),
    .io_s(HalfAdder_4_io_s),
    .io_co(HalfAdder_4_io_co)
  );
  HalfAdder HalfAdder_5 ( // @[wallace.scala 54:25]
    .io_a(HalfAdder_5_io_a),
    .io_b(HalfAdder_5_io_b),
    .io_s(HalfAdder_5_io_s),
    .io_co(HalfAdder_5_io_co)
  );
  FullAdder FullAdder_201 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_201_io_a),
    .io_b(FullAdder_201_io_b),
    .io_ci(FullAdder_201_io_ci),
    .io_s(FullAdder_201_io_s),
    .io_co(FullAdder_201_io_co)
  );
  FullAdder FullAdder_202 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_202_io_a),
    .io_b(FullAdder_202_io_b),
    .io_ci(FullAdder_202_io_ci),
    .io_s(FullAdder_202_io_s),
    .io_co(FullAdder_202_io_co)
  );
  FullAdder FullAdder_203 ( // @[wallace.scala 63:25]
    .io_a(FullAdder_203_io_a),
    .io_b(FullAdder_203_io_b),
    .io_ci(FullAdder_203_io_ci),
    .io_s(FullAdder_203_io_s),
    .io_co(FullAdder_203_io_co)
  );
  assign io_augend = {{1'd0}, _T_285}; // @[wallace.scala 86:13]
  assign io_addend = {{1'd0}, _T_315}; // @[wallace.scala 87:13]
  assign FullAdder_io_a = io_pp_13[15]; // @[wallace.scala 65:18]
  assign FullAdder_io_b = io_pp_14[14]; // @[wallace.scala 66:18]
  assign FullAdder_io_ci = io_pp_15[13]; // @[wallace.scala 67:19]
  assign FullAdder_1_io_a = io_pp_12[15]; // @[wallace.scala 65:18]
  assign FullAdder_1_io_b = io_pp_13[14]; // @[wallace.scala 66:18]
  assign FullAdder_1_io_ci = io_pp_14[13]; // @[wallace.scala 67:19]
  assign FullAdder_2_io_a = io_pp_11[15]; // @[wallace.scala 65:18]
  assign FullAdder_2_io_b = io_pp_12[14]; // @[wallace.scala 66:18]
  assign FullAdder_2_io_ci = io_pp_13[13]; // @[wallace.scala 67:19]
  assign FullAdder_3_io_a = io_pp_10[15]; // @[wallace.scala 65:18]
  assign FullAdder_3_io_b = io_pp_11[14]; // @[wallace.scala 66:18]
  assign FullAdder_3_io_ci = io_pp_12[13]; // @[wallace.scala 67:19]
  assign FullAdder_4_io_a = io_pp_13[12]; // @[wallace.scala 65:18]
  assign FullAdder_4_io_b = io_pp_14[11]; // @[wallace.scala 66:18]
  assign FullAdder_4_io_ci = io_pp_15[10]; // @[wallace.scala 67:19]
  assign FullAdder_5_io_a = io_pp_9[15]; // @[wallace.scala 65:18]
  assign FullAdder_5_io_b = io_pp_10[14]; // @[wallace.scala 66:18]
  assign FullAdder_5_io_ci = io_pp_11[13]; // @[wallace.scala 67:19]
  assign FullAdder_6_io_a = io_pp_12[12]; // @[wallace.scala 65:18]
  assign FullAdder_6_io_b = io_pp_13[11]; // @[wallace.scala 66:18]
  assign FullAdder_6_io_ci = io_pp_14[10]; // @[wallace.scala 67:19]
  assign FullAdder_7_io_a = io_pp_8[15]; // @[wallace.scala 65:18]
  assign FullAdder_7_io_b = io_pp_9[14]; // @[wallace.scala 66:18]
  assign FullAdder_7_io_ci = io_pp_10[13]; // @[wallace.scala 67:19]
  assign FullAdder_8_io_a = io_pp_11[12]; // @[wallace.scala 65:18]
  assign FullAdder_8_io_b = io_pp_12[11]; // @[wallace.scala 66:18]
  assign FullAdder_8_io_ci = io_pp_13[10]; // @[wallace.scala 67:19]
  assign FullAdder_9_io_a = io_pp_7[15]; // @[wallace.scala 65:18]
  assign FullAdder_9_io_b = io_pp_8[14]; // @[wallace.scala 66:18]
  assign FullAdder_9_io_ci = io_pp_9[13]; // @[wallace.scala 67:19]
  assign FullAdder_10_io_a = io_pp_10[12]; // @[wallace.scala 65:18]
  assign FullAdder_10_io_b = io_pp_11[11]; // @[wallace.scala 66:18]
  assign FullAdder_10_io_ci = io_pp_12[10]; // @[wallace.scala 67:19]
  assign FullAdder_11_io_a = io_pp_13[9]; // @[wallace.scala 65:18]
  assign FullAdder_11_io_b = io_pp_14[8]; // @[wallace.scala 66:18]
  assign FullAdder_11_io_ci = io_pp_15[7]; // @[wallace.scala 67:19]
  assign FullAdder_12_io_a = io_pp_6[15]; // @[wallace.scala 65:18]
  assign FullAdder_12_io_b = io_pp_7[14]; // @[wallace.scala 66:18]
  assign FullAdder_12_io_ci = io_pp_8[13]; // @[wallace.scala 67:19]
  assign FullAdder_13_io_a = io_pp_9[12]; // @[wallace.scala 65:18]
  assign FullAdder_13_io_b = io_pp_10[11]; // @[wallace.scala 66:18]
  assign FullAdder_13_io_ci = io_pp_11[10]; // @[wallace.scala 67:19]
  assign FullAdder_14_io_a = io_pp_12[9]; // @[wallace.scala 65:18]
  assign FullAdder_14_io_b = io_pp_13[8]; // @[wallace.scala 66:18]
  assign FullAdder_14_io_ci = io_pp_14[7]; // @[wallace.scala 67:19]
  assign FullAdder_15_io_a = io_pp_5[15]; // @[wallace.scala 65:18]
  assign FullAdder_15_io_b = io_pp_6[14]; // @[wallace.scala 66:18]
  assign FullAdder_15_io_ci = io_pp_7[13]; // @[wallace.scala 67:19]
  assign FullAdder_16_io_a = io_pp_8[12]; // @[wallace.scala 65:18]
  assign FullAdder_16_io_b = io_pp_9[11]; // @[wallace.scala 66:18]
  assign FullAdder_16_io_ci = io_pp_10[10]; // @[wallace.scala 67:19]
  assign FullAdder_17_io_a = io_pp_11[9]; // @[wallace.scala 65:18]
  assign FullAdder_17_io_b = io_pp_12[8]; // @[wallace.scala 66:18]
  assign FullAdder_17_io_ci = io_pp_13[7]; // @[wallace.scala 67:19]
  assign FullAdder_18_io_a = io_pp_4[15]; // @[wallace.scala 65:18]
  assign FullAdder_18_io_b = io_pp_5[14]; // @[wallace.scala 66:18]
  assign FullAdder_18_io_ci = io_pp_6[13]; // @[wallace.scala 67:19]
  assign FullAdder_19_io_a = io_pp_7[12]; // @[wallace.scala 65:18]
  assign FullAdder_19_io_b = io_pp_8[11]; // @[wallace.scala 66:18]
  assign FullAdder_19_io_ci = io_pp_9[10]; // @[wallace.scala 67:19]
  assign FullAdder_20_io_a = io_pp_10[9]; // @[wallace.scala 65:18]
  assign FullAdder_20_io_b = io_pp_11[8]; // @[wallace.scala 66:18]
  assign FullAdder_20_io_ci = io_pp_12[7]; // @[wallace.scala 67:19]
  assign FullAdder_21_io_a = io_pp_13[6]; // @[wallace.scala 65:18]
  assign FullAdder_21_io_b = io_pp_14[5]; // @[wallace.scala 66:18]
  assign FullAdder_21_io_ci = io_pp_15[4]; // @[wallace.scala 67:19]
  assign FullAdder_22_io_a = io_pp_3[15]; // @[wallace.scala 65:18]
  assign FullAdder_22_io_b = io_pp_4[14]; // @[wallace.scala 66:18]
  assign FullAdder_22_io_ci = io_pp_5[13]; // @[wallace.scala 67:19]
  assign FullAdder_23_io_a = io_pp_6[12]; // @[wallace.scala 65:18]
  assign FullAdder_23_io_b = io_pp_7[11]; // @[wallace.scala 66:18]
  assign FullAdder_23_io_ci = io_pp_8[10]; // @[wallace.scala 67:19]
  assign FullAdder_24_io_a = io_pp_9[9]; // @[wallace.scala 65:18]
  assign FullAdder_24_io_b = io_pp_10[8]; // @[wallace.scala 66:18]
  assign FullAdder_24_io_ci = io_pp_11[7]; // @[wallace.scala 67:19]
  assign FullAdder_25_io_a = io_pp_12[6]; // @[wallace.scala 65:18]
  assign FullAdder_25_io_b = io_pp_13[5]; // @[wallace.scala 66:18]
  assign FullAdder_25_io_ci = io_pp_14[4]; // @[wallace.scala 67:19]
  assign FullAdder_26_io_a = io_pp_2[15]; // @[wallace.scala 65:18]
  assign FullAdder_26_io_b = io_pp_3[14]; // @[wallace.scala 66:18]
  assign FullAdder_26_io_ci = io_pp_4[13]; // @[wallace.scala 67:19]
  assign FullAdder_27_io_a = io_pp_5[12]; // @[wallace.scala 65:18]
  assign FullAdder_27_io_b = io_pp_6[11]; // @[wallace.scala 66:18]
  assign FullAdder_27_io_ci = io_pp_7[10]; // @[wallace.scala 67:19]
  assign FullAdder_28_io_a = io_pp_8[9]; // @[wallace.scala 65:18]
  assign FullAdder_28_io_b = io_pp_9[8]; // @[wallace.scala 66:18]
  assign FullAdder_28_io_ci = io_pp_10[7]; // @[wallace.scala 67:19]
  assign FullAdder_29_io_a = io_pp_11[6]; // @[wallace.scala 65:18]
  assign FullAdder_29_io_b = io_pp_12[5]; // @[wallace.scala 66:18]
  assign FullAdder_29_io_ci = io_pp_13[4]; // @[wallace.scala 67:19]
  assign FullAdder_30_io_a = io_pp_1[15]; // @[wallace.scala 65:18]
  assign FullAdder_30_io_b = io_pp_2[14]; // @[wallace.scala 66:18]
  assign FullAdder_30_io_ci = io_pp_3[13]; // @[wallace.scala 67:19]
  assign FullAdder_31_io_a = io_pp_4[12]; // @[wallace.scala 65:18]
  assign FullAdder_31_io_b = io_pp_5[11]; // @[wallace.scala 66:18]
  assign FullAdder_31_io_ci = io_pp_6[10]; // @[wallace.scala 67:19]
  assign FullAdder_32_io_a = io_pp_7[9]; // @[wallace.scala 65:18]
  assign FullAdder_32_io_b = io_pp_8[8]; // @[wallace.scala 66:18]
  assign FullAdder_32_io_ci = io_pp_9[7]; // @[wallace.scala 67:19]
  assign FullAdder_33_io_a = io_pp_10[6]; // @[wallace.scala 65:18]
  assign FullAdder_33_io_b = io_pp_11[5]; // @[wallace.scala 66:18]
  assign FullAdder_33_io_ci = io_pp_12[4]; // @[wallace.scala 67:19]
  assign FullAdder_34_io_a = io_pp_13[3]; // @[wallace.scala 65:18]
  assign FullAdder_34_io_b = io_pp_14[2]; // @[wallace.scala 66:18]
  assign FullAdder_34_io_ci = io_pp_15[1]; // @[wallace.scala 67:19]
  assign FullAdder_35_io_a = io_pp_0[15]; // @[wallace.scala 65:18]
  assign FullAdder_35_io_b = io_pp_1[14]; // @[wallace.scala 66:18]
  assign FullAdder_35_io_ci = io_pp_2[13]; // @[wallace.scala 67:19]
  assign FullAdder_36_io_a = io_pp_3[12]; // @[wallace.scala 65:18]
  assign FullAdder_36_io_b = io_pp_4[11]; // @[wallace.scala 66:18]
  assign FullAdder_36_io_ci = io_pp_5[10]; // @[wallace.scala 67:19]
  assign FullAdder_37_io_a = io_pp_6[9]; // @[wallace.scala 65:18]
  assign FullAdder_37_io_b = io_pp_7[8]; // @[wallace.scala 66:18]
  assign FullAdder_37_io_ci = io_pp_8[7]; // @[wallace.scala 67:19]
  assign FullAdder_38_io_a = io_pp_9[6]; // @[wallace.scala 65:18]
  assign FullAdder_38_io_b = io_pp_10[5]; // @[wallace.scala 66:18]
  assign FullAdder_38_io_ci = io_pp_11[4]; // @[wallace.scala 67:19]
  assign FullAdder_39_io_a = io_pp_12[3]; // @[wallace.scala 65:18]
  assign FullAdder_39_io_b = io_pp_13[2]; // @[wallace.scala 66:18]
  assign FullAdder_39_io_ci = io_pp_14[1]; // @[wallace.scala 67:19]
  assign FullAdder_40_io_a = io_pp_0[14]; // @[wallace.scala 65:18]
  assign FullAdder_40_io_b = io_pp_1[13]; // @[wallace.scala 66:18]
  assign FullAdder_40_io_ci = io_pp_2[12]; // @[wallace.scala 67:19]
  assign FullAdder_41_io_a = io_pp_3[11]; // @[wallace.scala 65:18]
  assign FullAdder_41_io_b = io_pp_4[10]; // @[wallace.scala 66:18]
  assign FullAdder_41_io_ci = io_pp_5[9]; // @[wallace.scala 67:19]
  assign FullAdder_42_io_a = io_pp_6[8]; // @[wallace.scala 65:18]
  assign FullAdder_42_io_b = io_pp_7[7]; // @[wallace.scala 66:18]
  assign FullAdder_42_io_ci = io_pp_8[6]; // @[wallace.scala 67:19]
  assign FullAdder_43_io_a = io_pp_9[5]; // @[wallace.scala 65:18]
  assign FullAdder_43_io_b = io_pp_10[4]; // @[wallace.scala 66:18]
  assign FullAdder_43_io_ci = io_pp_11[3]; // @[wallace.scala 67:19]
  assign FullAdder_44_io_a = io_pp_12[2]; // @[wallace.scala 65:18]
  assign FullAdder_44_io_b = io_pp_13[1]; // @[wallace.scala 66:18]
  assign FullAdder_44_io_ci = io_pp_14[0]; // @[wallace.scala 67:19]
  assign FullAdder_45_io_a = io_pp_0[13]; // @[wallace.scala 65:18]
  assign FullAdder_45_io_b = io_pp_1[12]; // @[wallace.scala 66:18]
  assign FullAdder_45_io_ci = io_pp_2[11]; // @[wallace.scala 67:19]
  assign FullAdder_46_io_a = io_pp_3[10]; // @[wallace.scala 65:18]
  assign FullAdder_46_io_b = io_pp_4[9]; // @[wallace.scala 66:18]
  assign FullAdder_46_io_ci = io_pp_5[8]; // @[wallace.scala 67:19]
  assign FullAdder_47_io_a = io_pp_6[7]; // @[wallace.scala 65:18]
  assign FullAdder_47_io_b = io_pp_7[6]; // @[wallace.scala 66:18]
  assign FullAdder_47_io_ci = io_pp_8[5]; // @[wallace.scala 67:19]
  assign FullAdder_48_io_a = io_pp_9[4]; // @[wallace.scala 65:18]
  assign FullAdder_48_io_b = io_pp_10[3]; // @[wallace.scala 66:18]
  assign FullAdder_48_io_ci = io_pp_11[2]; // @[wallace.scala 67:19]
  assign FullAdder_49_io_a = io_pp_0[12]; // @[wallace.scala 65:18]
  assign FullAdder_49_io_b = io_pp_1[11]; // @[wallace.scala 66:18]
  assign FullAdder_49_io_ci = io_pp_2[10]; // @[wallace.scala 67:19]
  assign FullAdder_50_io_a = io_pp_3[9]; // @[wallace.scala 65:18]
  assign FullAdder_50_io_b = io_pp_4[8]; // @[wallace.scala 66:18]
  assign FullAdder_50_io_ci = io_pp_5[7]; // @[wallace.scala 67:19]
  assign FullAdder_51_io_a = io_pp_6[6]; // @[wallace.scala 65:18]
  assign FullAdder_51_io_b = io_pp_7[5]; // @[wallace.scala 66:18]
  assign FullAdder_51_io_ci = io_pp_8[4]; // @[wallace.scala 67:19]
  assign FullAdder_52_io_a = io_pp_9[3]; // @[wallace.scala 65:18]
  assign FullAdder_52_io_b = io_pp_10[2]; // @[wallace.scala 66:18]
  assign FullAdder_52_io_ci = io_pp_11[1]; // @[wallace.scala 67:19]
  assign FullAdder_53_io_a = io_pp_0[11]; // @[wallace.scala 65:18]
  assign FullAdder_53_io_b = io_pp_1[10]; // @[wallace.scala 66:18]
  assign FullAdder_53_io_ci = io_pp_2[9]; // @[wallace.scala 67:19]
  assign FullAdder_54_io_a = io_pp_3[8]; // @[wallace.scala 65:18]
  assign FullAdder_54_io_b = io_pp_4[7]; // @[wallace.scala 66:18]
  assign FullAdder_54_io_ci = io_pp_5[6]; // @[wallace.scala 67:19]
  assign FullAdder_55_io_a = io_pp_6[5]; // @[wallace.scala 65:18]
  assign FullAdder_55_io_b = io_pp_7[4]; // @[wallace.scala 66:18]
  assign FullAdder_55_io_ci = io_pp_8[3]; // @[wallace.scala 67:19]
  assign FullAdder_56_io_a = io_pp_9[2]; // @[wallace.scala 65:18]
  assign FullAdder_56_io_b = io_pp_10[1]; // @[wallace.scala 66:18]
  assign FullAdder_56_io_ci = io_pp_11[0]; // @[wallace.scala 67:19]
  assign FullAdder_57_io_a = io_pp_0[10]; // @[wallace.scala 65:18]
  assign FullAdder_57_io_b = io_pp_1[9]; // @[wallace.scala 66:18]
  assign FullAdder_57_io_ci = io_pp_2[8]; // @[wallace.scala 67:19]
  assign FullAdder_58_io_a = io_pp_3[7]; // @[wallace.scala 65:18]
  assign FullAdder_58_io_b = io_pp_4[6]; // @[wallace.scala 66:18]
  assign FullAdder_58_io_ci = io_pp_5[5]; // @[wallace.scala 67:19]
  assign FullAdder_59_io_a = io_pp_6[4]; // @[wallace.scala 65:18]
  assign FullAdder_59_io_b = io_pp_7[3]; // @[wallace.scala 66:18]
  assign FullAdder_59_io_ci = io_pp_8[2]; // @[wallace.scala 67:19]
  assign FullAdder_60_io_a = io_pp_0[9]; // @[wallace.scala 65:18]
  assign FullAdder_60_io_b = io_pp_1[8]; // @[wallace.scala 66:18]
  assign FullAdder_60_io_ci = io_pp_2[7]; // @[wallace.scala 67:19]
  assign FullAdder_61_io_a = io_pp_3[6]; // @[wallace.scala 65:18]
  assign FullAdder_61_io_b = io_pp_4[5]; // @[wallace.scala 66:18]
  assign FullAdder_61_io_ci = io_pp_5[4]; // @[wallace.scala 67:19]
  assign FullAdder_62_io_a = io_pp_6[3]; // @[wallace.scala 65:18]
  assign FullAdder_62_io_b = io_pp_7[2]; // @[wallace.scala 66:18]
  assign FullAdder_62_io_ci = io_pp_8[1]; // @[wallace.scala 67:19]
  assign FullAdder_63_io_a = io_pp_0[8]; // @[wallace.scala 65:18]
  assign FullAdder_63_io_b = io_pp_1[7]; // @[wallace.scala 66:18]
  assign FullAdder_63_io_ci = io_pp_2[6]; // @[wallace.scala 67:19]
  assign FullAdder_64_io_a = io_pp_3[5]; // @[wallace.scala 65:18]
  assign FullAdder_64_io_b = io_pp_4[4]; // @[wallace.scala 66:18]
  assign FullAdder_64_io_ci = io_pp_5[3]; // @[wallace.scala 67:19]
  assign FullAdder_65_io_a = io_pp_6[2]; // @[wallace.scala 65:18]
  assign FullAdder_65_io_b = io_pp_7[1]; // @[wallace.scala 66:18]
  assign FullAdder_65_io_ci = io_pp_8[0]; // @[wallace.scala 67:19]
  assign FullAdder_66_io_a = io_pp_0[7]; // @[wallace.scala 65:18]
  assign FullAdder_66_io_b = io_pp_1[6]; // @[wallace.scala 66:18]
  assign FullAdder_66_io_ci = io_pp_2[5]; // @[wallace.scala 67:19]
  assign FullAdder_67_io_a = io_pp_3[4]; // @[wallace.scala 65:18]
  assign FullAdder_67_io_b = io_pp_4[3]; // @[wallace.scala 66:18]
  assign FullAdder_67_io_ci = io_pp_5[2]; // @[wallace.scala 67:19]
  assign FullAdder_68_io_a = io_pp_0[6]; // @[wallace.scala 65:18]
  assign FullAdder_68_io_b = io_pp_1[5]; // @[wallace.scala 66:18]
  assign FullAdder_68_io_ci = io_pp_2[4]; // @[wallace.scala 67:19]
  assign FullAdder_69_io_a = io_pp_3[3]; // @[wallace.scala 65:18]
  assign FullAdder_69_io_b = io_pp_4[2]; // @[wallace.scala 66:18]
  assign FullAdder_69_io_ci = io_pp_5[1]; // @[wallace.scala 67:19]
  assign FullAdder_70_io_a = io_pp_0[5]; // @[wallace.scala 65:18]
  assign FullAdder_70_io_b = io_pp_1[4]; // @[wallace.scala 66:18]
  assign FullAdder_70_io_ci = io_pp_2[3]; // @[wallace.scala 67:19]
  assign FullAdder_71_io_a = io_pp_3[2]; // @[wallace.scala 65:18]
  assign FullAdder_71_io_b = io_pp_4[1]; // @[wallace.scala 66:18]
  assign FullAdder_71_io_ci = io_pp_5[0]; // @[wallace.scala 67:19]
  assign FullAdder_72_io_a = io_pp_0[4]; // @[wallace.scala 65:18]
  assign FullAdder_72_io_b = io_pp_1[3]; // @[wallace.scala 66:18]
  assign FullAdder_72_io_ci = io_pp_2[2]; // @[wallace.scala 67:19]
  assign FullAdder_73_io_a = io_pp_0[3]; // @[wallace.scala 65:18]
  assign FullAdder_73_io_b = io_pp_1[2]; // @[wallace.scala 66:18]
  assign FullAdder_73_io_ci = io_pp_2[1]; // @[wallace.scala 67:19]
  assign FullAdder_74_io_a = io_pp_0[2]; // @[wallace.scala 65:18]
  assign FullAdder_74_io_b = io_pp_1[1]; // @[wallace.scala 66:18]
  assign FullAdder_74_io_ci = io_pp_2[0]; // @[wallace.scala 67:19]
  assign FullAdder_75_io_a = io_pp_14[15]; // @[wallace.scala 65:18]
  assign FullAdder_75_io_b = io_pp_15[14]; // @[wallace.scala 66:18]
  assign FullAdder_75_io_ci = FullAdder_io_co; // @[wallace.scala 67:19]
  assign FullAdder_76_io_a = io_pp_15[12]; // @[wallace.scala 65:18]
  assign FullAdder_76_io_b = FullAdder_1_io_s; // @[wallace.scala 66:18]
  assign FullAdder_76_io_ci = FullAdder_2_io_co; // @[wallace.scala 67:19]
  assign FullAdder_77_io_a = io_pp_14[12]; // @[wallace.scala 65:18]
  assign FullAdder_77_io_b = io_pp_15[11]; // @[wallace.scala 66:18]
  assign FullAdder_77_io_ci = FullAdder_2_io_s; // @[wallace.scala 67:19]
  assign FullAdder_78_io_a = FullAdder_3_io_s; // @[wallace.scala 65:18]
  assign FullAdder_78_io_b = FullAdder_4_io_s; // @[wallace.scala 66:18]
  assign FullAdder_78_io_ci = FullAdder_5_io_co; // @[wallace.scala 67:19]
  assign FullAdder_79_io_a = io_pp_15[9]; // @[wallace.scala 65:18]
  assign FullAdder_79_io_b = FullAdder_5_io_s; // @[wallace.scala 66:18]
  assign FullAdder_79_io_ci = FullAdder_6_io_s; // @[wallace.scala 67:19]
  assign FullAdder_80_io_a = io_pp_14[9]; // @[wallace.scala 65:18]
  assign FullAdder_80_io_b = io_pp_15[8]; // @[wallace.scala 66:18]
  assign FullAdder_80_io_ci = FullAdder_7_io_s; // @[wallace.scala 67:19]
  assign FullAdder_81_io_a = FullAdder_8_io_s; // @[wallace.scala 65:18]
  assign FullAdder_81_io_b = FullAdder_9_io_co; // @[wallace.scala 66:18]
  assign FullAdder_81_io_ci = FullAdder_10_io_co; // @[wallace.scala 67:19]
  assign FullAdder_82_io_a = FullAdder_9_io_s; // @[wallace.scala 65:18]
  assign FullAdder_82_io_b = FullAdder_10_io_s; // @[wallace.scala 66:18]
  assign FullAdder_82_io_ci = FullAdder_11_io_s; // @[wallace.scala 67:19]
  assign FullAdder_83_io_a = FullAdder_12_io_co; // @[wallace.scala 65:18]
  assign FullAdder_83_io_b = FullAdder_13_io_co; // @[wallace.scala 66:18]
  assign FullAdder_83_io_ci = FullAdder_14_io_co; // @[wallace.scala 67:19]
  assign FullAdder_84_io_a = io_pp_15[6]; // @[wallace.scala 65:18]
  assign FullAdder_84_io_b = FullAdder_12_io_s; // @[wallace.scala 66:18]
  assign FullAdder_84_io_ci = FullAdder_13_io_s; // @[wallace.scala 67:19]
  assign FullAdder_85_io_a = FullAdder_14_io_s; // @[wallace.scala 65:18]
  assign FullAdder_85_io_b = FullAdder_15_io_co; // @[wallace.scala 66:18]
  assign FullAdder_85_io_ci = FullAdder_16_io_co; // @[wallace.scala 67:19]
  assign FullAdder_86_io_a = io_pp_14[6]; // @[wallace.scala 65:18]
  assign FullAdder_86_io_b = io_pp_15[5]; // @[wallace.scala 66:18]
  assign FullAdder_86_io_ci = FullAdder_15_io_s; // @[wallace.scala 67:19]
  assign FullAdder_87_io_a = FullAdder_16_io_s; // @[wallace.scala 65:18]
  assign FullAdder_87_io_b = FullAdder_17_io_s; // @[wallace.scala 66:18]
  assign FullAdder_87_io_ci = FullAdder_18_io_co; // @[wallace.scala 67:19]
  assign FullAdder_88_io_a = FullAdder_19_io_co; // @[wallace.scala 65:18]
  assign FullAdder_88_io_b = FullAdder_20_io_co; // @[wallace.scala 66:18]
  assign FullAdder_88_io_ci = FullAdder_21_io_co; // @[wallace.scala 67:19]
  assign FullAdder_89_io_a = FullAdder_18_io_s; // @[wallace.scala 65:18]
  assign FullAdder_89_io_b = FullAdder_19_io_s; // @[wallace.scala 66:18]
  assign FullAdder_89_io_ci = FullAdder_20_io_s; // @[wallace.scala 67:19]
  assign FullAdder_90_io_a = FullAdder_21_io_s; // @[wallace.scala 65:18]
  assign FullAdder_90_io_b = FullAdder_22_io_co; // @[wallace.scala 66:18]
  assign FullAdder_90_io_ci = FullAdder_23_io_co; // @[wallace.scala 67:19]
  assign FullAdder_91_io_a = io_pp_15[3]; // @[wallace.scala 65:18]
  assign FullAdder_91_io_b = FullAdder_22_io_s; // @[wallace.scala 66:18]
  assign FullAdder_91_io_ci = FullAdder_23_io_s; // @[wallace.scala 67:19]
  assign FullAdder_92_io_a = FullAdder_24_io_s; // @[wallace.scala 65:18]
  assign FullAdder_92_io_b = FullAdder_25_io_s; // @[wallace.scala 66:18]
  assign FullAdder_92_io_ci = FullAdder_26_io_co; // @[wallace.scala 67:19]
  assign FullAdder_93_io_a = FullAdder_27_io_co; // @[wallace.scala 65:18]
  assign FullAdder_93_io_b = FullAdder_28_io_co; // @[wallace.scala 66:18]
  assign FullAdder_93_io_ci = FullAdder_29_io_co; // @[wallace.scala 67:19]
  assign FullAdder_94_io_a = io_pp_14[3]; // @[wallace.scala 65:18]
  assign FullAdder_94_io_b = io_pp_15[2]; // @[wallace.scala 66:18]
  assign FullAdder_94_io_ci = FullAdder_26_io_s; // @[wallace.scala 67:19]
  assign FullAdder_95_io_a = FullAdder_27_io_s; // @[wallace.scala 65:18]
  assign FullAdder_95_io_b = FullAdder_28_io_s; // @[wallace.scala 66:18]
  assign FullAdder_95_io_ci = FullAdder_29_io_s; // @[wallace.scala 67:19]
  assign FullAdder_96_io_a = FullAdder_30_io_co; // @[wallace.scala 65:18]
  assign FullAdder_96_io_b = FullAdder_31_io_co; // @[wallace.scala 66:18]
  assign FullAdder_96_io_ci = FullAdder_32_io_co; // @[wallace.scala 67:19]
  assign FullAdder_97_io_a = FullAdder_30_io_s; // @[wallace.scala 65:18]
  assign FullAdder_97_io_b = FullAdder_31_io_s; // @[wallace.scala 66:18]
  assign FullAdder_97_io_ci = FullAdder_32_io_s; // @[wallace.scala 67:19]
  assign FullAdder_98_io_a = FullAdder_33_io_s; // @[wallace.scala 65:18]
  assign FullAdder_98_io_b = FullAdder_34_io_s; // @[wallace.scala 66:18]
  assign FullAdder_98_io_ci = FullAdder_35_io_co; // @[wallace.scala 67:19]
  assign FullAdder_99_io_a = FullAdder_36_io_co; // @[wallace.scala 65:18]
  assign FullAdder_99_io_b = FullAdder_37_io_co; // @[wallace.scala 66:18]
  assign FullAdder_99_io_ci = FullAdder_38_io_co; // @[wallace.scala 67:19]
  assign FullAdder_100_io_a = io_pp_15[0]; // @[wallace.scala 65:18]
  assign FullAdder_100_io_b = FullAdder_35_io_s; // @[wallace.scala 66:18]
  assign FullAdder_100_io_ci = FullAdder_36_io_s; // @[wallace.scala 67:19]
  assign FullAdder_101_io_a = FullAdder_37_io_s; // @[wallace.scala 65:18]
  assign FullAdder_101_io_b = FullAdder_38_io_s; // @[wallace.scala 66:18]
  assign FullAdder_101_io_ci = FullAdder_39_io_s; // @[wallace.scala 67:19]
  assign FullAdder_102_io_a = FullAdder_40_io_co; // @[wallace.scala 65:18]
  assign FullAdder_102_io_b = FullAdder_41_io_co; // @[wallace.scala 66:18]
  assign FullAdder_102_io_ci = FullAdder_42_io_co; // @[wallace.scala 67:19]
  assign FullAdder_103_io_a = FullAdder_40_io_s; // @[wallace.scala 65:18]
  assign FullAdder_103_io_b = FullAdder_41_io_s; // @[wallace.scala 66:18]
  assign FullAdder_103_io_ci = FullAdder_42_io_s; // @[wallace.scala 67:19]
  assign FullAdder_104_io_a = FullAdder_43_io_s; // @[wallace.scala 65:18]
  assign FullAdder_104_io_b = FullAdder_44_io_s; // @[wallace.scala 66:18]
  assign FullAdder_104_io_ci = FullAdder_45_io_co; // @[wallace.scala 67:19]
  assign FullAdder_105_io_a = FullAdder_46_io_co; // @[wallace.scala 65:18]
  assign FullAdder_105_io_b = FullAdder_47_io_co; // @[wallace.scala 66:18]
  assign FullAdder_105_io_ci = FullAdder_48_io_co; // @[wallace.scala 67:19]
  assign FullAdder_106_io_a = io_pp_12[1]; // @[wallace.scala 65:18]
  assign FullAdder_106_io_b = io_pp_13[0]; // @[wallace.scala 66:18]
  assign FullAdder_106_io_ci = FullAdder_45_io_s; // @[wallace.scala 67:19]
  assign FullAdder_107_io_a = FullAdder_46_io_s; // @[wallace.scala 65:18]
  assign FullAdder_107_io_b = FullAdder_47_io_s; // @[wallace.scala 66:18]
  assign FullAdder_107_io_ci = FullAdder_48_io_s; // @[wallace.scala 67:19]
  assign FullAdder_108_io_a = FullAdder_49_io_co; // @[wallace.scala 65:18]
  assign FullAdder_108_io_b = FullAdder_50_io_co; // @[wallace.scala 66:18]
  assign FullAdder_108_io_ci = FullAdder_51_io_co; // @[wallace.scala 67:19]
  assign FullAdder_109_io_a = io_pp_12[0]; // @[wallace.scala 65:18]
  assign FullAdder_109_io_b = FullAdder_49_io_s; // @[wallace.scala 66:18]
  assign FullAdder_109_io_ci = FullAdder_50_io_s; // @[wallace.scala 67:19]
  assign FullAdder_110_io_a = FullAdder_51_io_s; // @[wallace.scala 65:18]
  assign FullAdder_110_io_b = FullAdder_52_io_s; // @[wallace.scala 66:18]
  assign FullAdder_110_io_ci = FullAdder_53_io_co; // @[wallace.scala 67:19]
  assign FullAdder_111_io_a = FullAdder_54_io_co; // @[wallace.scala 65:18]
  assign FullAdder_111_io_b = FullAdder_55_io_co; // @[wallace.scala 66:18]
  assign FullAdder_111_io_ci = FullAdder_56_io_co; // @[wallace.scala 67:19]
  assign FullAdder_112_io_a = FullAdder_53_io_s; // @[wallace.scala 65:18]
  assign FullAdder_112_io_b = FullAdder_54_io_s; // @[wallace.scala 66:18]
  assign FullAdder_112_io_ci = FullAdder_55_io_s; // @[wallace.scala 67:19]
  assign FullAdder_113_io_a = FullAdder_56_io_s; // @[wallace.scala 65:18]
  assign FullAdder_113_io_b = FullAdder_57_io_co; // @[wallace.scala 66:18]
  assign FullAdder_113_io_ci = FullAdder_58_io_co; // @[wallace.scala 67:19]
  assign FullAdder_114_io_a = io_pp_9[1]; // @[wallace.scala 65:18]
  assign FullAdder_114_io_b = io_pp_10[0]; // @[wallace.scala 66:18]
  assign FullAdder_114_io_ci = FullAdder_57_io_s; // @[wallace.scala 67:19]
  assign FullAdder_115_io_a = FullAdder_58_io_s; // @[wallace.scala 65:18]
  assign FullAdder_115_io_b = FullAdder_59_io_s; // @[wallace.scala 66:18]
  assign FullAdder_115_io_ci = FullAdder_60_io_co; // @[wallace.scala 67:19]
  assign FullAdder_116_io_a = io_pp_9[0]; // @[wallace.scala 65:18]
  assign FullAdder_116_io_b = FullAdder_60_io_s; // @[wallace.scala 66:18]
  assign FullAdder_116_io_ci = FullAdder_61_io_s; // @[wallace.scala 67:19]
  assign FullAdder_117_io_a = FullAdder_62_io_s; // @[wallace.scala 65:18]
  assign FullAdder_117_io_b = FullAdder_63_io_co; // @[wallace.scala 66:18]
  assign FullAdder_117_io_ci = FullAdder_64_io_co; // @[wallace.scala 67:19]
  assign FullAdder_118_io_a = FullAdder_63_io_s; // @[wallace.scala 65:18]
  assign FullAdder_118_io_b = FullAdder_64_io_s; // @[wallace.scala 66:18]
  assign FullAdder_118_io_ci = FullAdder_65_io_s; // @[wallace.scala 67:19]
  assign FullAdder_119_io_a = io_pp_6[1]; // @[wallace.scala 65:18]
  assign FullAdder_119_io_b = io_pp_7[0]; // @[wallace.scala 66:18]
  assign FullAdder_119_io_ci = FullAdder_66_io_s; // @[wallace.scala 67:19]
  assign FullAdder_120_io_a = FullAdder_67_io_s; // @[wallace.scala 65:18]
  assign FullAdder_120_io_b = FullAdder_68_io_co; // @[wallace.scala 66:18]
  assign FullAdder_120_io_ci = FullAdder_69_io_co; // @[wallace.scala 67:19]
  assign FullAdder_121_io_a = io_pp_6[0]; // @[wallace.scala 65:18]
  assign FullAdder_121_io_b = FullAdder_68_io_s; // @[wallace.scala 66:18]
  assign FullAdder_121_io_ci = FullAdder_69_io_s; // @[wallace.scala 67:19]
  assign FullAdder_122_io_a = FullAdder_70_io_s; // @[wallace.scala 65:18]
  assign FullAdder_122_io_b = FullAdder_71_io_s; // @[wallace.scala 66:18]
  assign FullAdder_122_io_ci = FullAdder_72_io_co; // @[wallace.scala 67:19]
  assign FullAdder_123_io_a = io_pp_3[1]; // @[wallace.scala 65:18]
  assign FullAdder_123_io_b = io_pp_4[0]; // @[wallace.scala 66:18]
  assign FullAdder_123_io_ci = FullAdder_72_io_s; // @[wallace.scala 67:19]
  assign FullAdder_124_io_a = io_pp_3[0]; // @[wallace.scala 65:18]
  assign FullAdder_124_io_b = FullAdder_73_io_s; // @[wallace.scala 66:18]
  assign FullAdder_124_io_ci = FullAdder_74_io_co; // @[wallace.scala 67:19]
  assign FullAdder_125_io_a = FullAdder_io_s; // @[wallace.scala 65:18]
  assign FullAdder_125_io_b = FullAdder_1_io_co; // @[wallace.scala 66:18]
  assign FullAdder_125_io_ci = FullAdder_76_io_co; // @[wallace.scala 67:19]
  assign FullAdder_126_io_a = FullAdder_3_io_co; // @[wallace.scala 65:18]
  assign FullAdder_126_io_b = FullAdder_4_io_co; // @[wallace.scala 66:18]
  assign FullAdder_126_io_ci = FullAdder_77_io_s; // @[wallace.scala 67:19]
  assign FullAdder_127_io_a = FullAdder_6_io_co; // @[wallace.scala 65:18]
  assign FullAdder_127_io_b = FullAdder_78_io_s; // @[wallace.scala 66:18]
  assign FullAdder_127_io_ci = FullAdder_79_io_co; // @[wallace.scala 67:19]
  assign FullAdder_128_io_a = FullAdder_7_io_co; // @[wallace.scala 65:18]
  assign FullAdder_128_io_b = FullAdder_8_io_co; // @[wallace.scala 66:18]
  assign FullAdder_128_io_ci = FullAdder_79_io_s; // @[wallace.scala 67:19]
  assign FullAdder_129_io_a = FullAdder_11_io_co; // @[wallace.scala 65:18]
  assign FullAdder_129_io_b = FullAdder_80_io_s; // @[wallace.scala 66:18]
  assign FullAdder_129_io_ci = FullAdder_81_io_s; // @[wallace.scala 67:19]
  assign FullAdder_130_io_a = FullAdder_82_io_s; // @[wallace.scala 65:18]
  assign FullAdder_130_io_b = FullAdder_83_io_s; // @[wallace.scala 66:18]
  assign FullAdder_130_io_ci = FullAdder_84_io_co; // @[wallace.scala 67:19]
  assign FullAdder_131_io_a = FullAdder_17_io_co; // @[wallace.scala 65:18]
  assign FullAdder_131_io_b = FullAdder_84_io_s; // @[wallace.scala 66:18]
  assign FullAdder_131_io_ci = FullAdder_85_io_s; // @[wallace.scala 67:19]
  assign FullAdder_132_io_a = FullAdder_86_io_co; // @[wallace.scala 65:18]
  assign FullAdder_132_io_b = FullAdder_87_io_co; // @[wallace.scala 66:18]
  assign FullAdder_132_io_ci = FullAdder_88_io_co; // @[wallace.scala 67:19]
  assign FullAdder_133_io_a = FullAdder_86_io_s; // @[wallace.scala 65:18]
  assign FullAdder_133_io_b = FullAdder_87_io_s; // @[wallace.scala 66:18]
  assign FullAdder_133_io_ci = FullAdder_88_io_s; // @[wallace.scala 67:19]
  assign FullAdder_134_io_a = FullAdder_24_io_co; // @[wallace.scala 65:18]
  assign FullAdder_134_io_b = FullAdder_25_io_co; // @[wallace.scala 66:18]
  assign FullAdder_134_io_ci = FullAdder_89_io_s; // @[wallace.scala 67:19]
  assign FullAdder_135_io_a = FullAdder_90_io_s; // @[wallace.scala 65:18]
  assign FullAdder_135_io_b = FullAdder_91_io_co; // @[wallace.scala 66:18]
  assign FullAdder_135_io_ci = FullAdder_92_io_co; // @[wallace.scala 67:19]
  assign FullAdder_136_io_a = FullAdder_91_io_s; // @[wallace.scala 65:18]
  assign FullAdder_136_io_b = FullAdder_92_io_s; // @[wallace.scala 66:18]
  assign FullAdder_136_io_ci = FullAdder_93_io_s; // @[wallace.scala 67:19]
  assign FullAdder_137_io_a = FullAdder_94_io_co; // @[wallace.scala 65:18]
  assign FullAdder_137_io_b = FullAdder_95_io_co; // @[wallace.scala 66:18]
  assign FullAdder_137_io_ci = FullAdder_96_io_co; // @[wallace.scala 67:19]
  assign FullAdder_138_io_a = FullAdder_33_io_co; // @[wallace.scala 65:18]
  assign FullAdder_138_io_b = FullAdder_34_io_co; // @[wallace.scala 66:18]
  assign FullAdder_138_io_ci = FullAdder_94_io_s; // @[wallace.scala 67:19]
  assign FullAdder_139_io_a = FullAdder_95_io_s; // @[wallace.scala 65:18]
  assign FullAdder_139_io_b = FullAdder_96_io_s; // @[wallace.scala 66:18]
  assign FullAdder_139_io_ci = FullAdder_97_io_co; // @[wallace.scala 67:19]
  assign FullAdder_140_io_a = FullAdder_39_io_co; // @[wallace.scala 65:18]
  assign FullAdder_140_io_b = FullAdder_97_io_s; // @[wallace.scala 66:18]
  assign FullAdder_140_io_ci = FullAdder_98_io_s; // @[wallace.scala 67:19]
  assign FullAdder_141_io_a = FullAdder_99_io_s; // @[wallace.scala 65:18]
  assign FullAdder_141_io_b = FullAdder_100_io_co; // @[wallace.scala 66:18]
  assign FullAdder_141_io_ci = FullAdder_101_io_co; // @[wallace.scala 67:19]
  assign FullAdder_142_io_a = FullAdder_43_io_co; // @[wallace.scala 65:18]
  assign FullAdder_142_io_b = FullAdder_44_io_co; // @[wallace.scala 66:18]
  assign FullAdder_142_io_ci = FullAdder_100_io_s; // @[wallace.scala 67:19]
  assign FullAdder_143_io_a = FullAdder_101_io_s; // @[wallace.scala 65:18]
  assign FullAdder_143_io_b = FullAdder_102_io_s; // @[wallace.scala 66:18]
  assign FullAdder_143_io_ci = FullAdder_103_io_co; // @[wallace.scala 67:19]
  assign FullAdder_144_io_a = FullAdder_103_io_s; // @[wallace.scala 65:18]
  assign FullAdder_144_io_b = FullAdder_104_io_s; // @[wallace.scala 66:18]
  assign FullAdder_144_io_ci = FullAdder_105_io_s; // @[wallace.scala 67:19]
  assign FullAdder_145_io_a = FullAdder_106_io_co; // @[wallace.scala 65:18]
  assign FullAdder_145_io_b = FullAdder_107_io_co; // @[wallace.scala 66:18]
  assign FullAdder_145_io_ci = FullAdder_108_io_co; // @[wallace.scala 67:19]
  assign FullAdder_146_io_a = FullAdder_52_io_co; // @[wallace.scala 65:18]
  assign FullAdder_146_io_b = FullAdder_106_io_s; // @[wallace.scala 66:18]
  assign FullAdder_146_io_ci = FullAdder_107_io_s; // @[wallace.scala 67:19]
  assign FullAdder_147_io_a = FullAdder_108_io_s; // @[wallace.scala 65:18]
  assign FullAdder_147_io_b = FullAdder_109_io_co; // @[wallace.scala 66:18]
  assign FullAdder_147_io_ci = FullAdder_110_io_co; // @[wallace.scala 67:19]
  assign FullAdder_148_io_a = FullAdder_109_io_s; // @[wallace.scala 65:18]
  assign FullAdder_148_io_b = FullAdder_110_io_s; // @[wallace.scala 66:18]
  assign FullAdder_148_io_ci = FullAdder_111_io_s; // @[wallace.scala 67:19]
  assign FullAdder_149_io_a = FullAdder_59_io_co; // @[wallace.scala 65:18]
  assign FullAdder_149_io_b = FullAdder_112_io_s; // @[wallace.scala 66:18]
  assign FullAdder_149_io_ci = FullAdder_113_io_s; // @[wallace.scala 67:19]
  assign FullAdder_150_io_a = FullAdder_61_io_co; // @[wallace.scala 65:18]
  assign FullAdder_150_io_b = FullAdder_62_io_co; // @[wallace.scala 66:18]
  assign FullAdder_150_io_ci = FullAdder_114_io_s; // @[wallace.scala 67:19]
  assign FullAdder_151_io_a = FullAdder_115_io_s; // @[wallace.scala 65:18]
  assign FullAdder_151_io_b = FullAdder_116_io_co; // @[wallace.scala 66:18]
  assign FullAdder_151_io_ci = FullAdder_117_io_co; // @[wallace.scala 67:19]
  assign FullAdder_152_io_a = FullAdder_65_io_co; // @[wallace.scala 65:18]
  assign FullAdder_152_io_b = FullAdder_116_io_s; // @[wallace.scala 66:18]
  assign FullAdder_152_io_ci = FullAdder_117_io_s; // @[wallace.scala 67:19]
  assign FullAdder_153_io_a = FullAdder_66_io_co; // @[wallace.scala 65:18]
  assign FullAdder_153_io_b = FullAdder_67_io_co; // @[wallace.scala 66:18]
  assign FullAdder_153_io_ci = FullAdder_118_io_s; // @[wallace.scala 67:19]
  assign HalfAdder_io_a = FullAdder_119_io_co; // @[wallace.scala 56:18]
  assign HalfAdder_io_b = FullAdder_120_io_co; // @[wallace.scala 57:18]
  assign FullAdder_154_io_a = FullAdder_119_io_s; // @[wallace.scala 65:18]
  assign FullAdder_154_io_b = FullAdder_120_io_s; // @[wallace.scala 66:18]
  assign FullAdder_154_io_ci = FullAdder_121_io_co; // @[wallace.scala 67:19]
  assign FullAdder_155_io_a = FullAdder_70_io_co; // @[wallace.scala 65:18]
  assign FullAdder_155_io_b = FullAdder_71_io_co; // @[wallace.scala 66:18]
  assign FullAdder_155_io_ci = FullAdder_121_io_s; // @[wallace.scala 67:19]
  assign FullAdder_156_io_a = FullAdder_73_io_co; // @[wallace.scala 65:18]
  assign FullAdder_156_io_b = FullAdder_123_io_s; // @[wallace.scala 66:18]
  assign FullAdder_156_io_ci = FullAdder_124_io_co; // @[wallace.scala 67:19]
  assign FullAdder_157_io_a = FullAdder_76_io_s; // @[wallace.scala 65:18]
  assign FullAdder_157_io_b = FullAdder_77_io_co; // @[wallace.scala 66:18]
  assign FullAdder_157_io_ci = FullAdder_126_io_co; // @[wallace.scala 67:19]
  assign FullAdder_158_io_a = FullAdder_78_io_co; // @[wallace.scala 65:18]
  assign FullAdder_158_io_b = FullAdder_126_io_s; // @[wallace.scala 66:18]
  assign FullAdder_158_io_ci = FullAdder_127_io_co; // @[wallace.scala 67:19]
  assign FullAdder_159_io_a = FullAdder_80_io_co; // @[wallace.scala 65:18]
  assign FullAdder_159_io_b = FullAdder_81_io_co; // @[wallace.scala 66:18]
  assign FullAdder_159_io_ci = FullAdder_128_io_s; // @[wallace.scala 67:19]
  assign FullAdder_160_io_a = FullAdder_82_io_co; // @[wallace.scala 65:18]
  assign FullAdder_160_io_b = FullAdder_83_io_co; // @[wallace.scala 66:18]
  assign FullAdder_160_io_ci = FullAdder_129_io_s; // @[wallace.scala 67:19]
  assign FullAdder_161_io_a = FullAdder_85_io_co; // @[wallace.scala 65:18]
  assign FullAdder_161_io_b = FullAdder_130_io_s; // @[wallace.scala 66:18]
  assign FullAdder_161_io_ci = FullAdder_131_io_co; // @[wallace.scala 67:19]
  assign FullAdder_162_io_a = FullAdder_131_io_s; // @[wallace.scala 65:18]
  assign FullAdder_162_io_b = FullAdder_132_io_s; // @[wallace.scala 66:18]
  assign FullAdder_162_io_ci = FullAdder_133_io_co; // @[wallace.scala 67:19]
  assign FullAdder_163_io_a = FullAdder_89_io_co; // @[wallace.scala 65:18]
  assign FullAdder_163_io_b = FullAdder_90_io_co; // @[wallace.scala 66:18]
  assign FullAdder_163_io_ci = FullAdder_133_io_s; // @[wallace.scala 67:19]
  assign FullAdder_164_io_a = FullAdder_93_io_co; // @[wallace.scala 65:18]
  assign FullAdder_164_io_b = FullAdder_134_io_s; // @[wallace.scala 66:18]
  assign FullAdder_164_io_ci = FullAdder_135_io_s; // @[wallace.scala 67:19]
  assign FullAdder_165_io_a = FullAdder_136_io_s; // @[wallace.scala 65:18]
  assign FullAdder_165_io_b = FullAdder_137_io_s; // @[wallace.scala 66:18]
  assign FullAdder_165_io_ci = FullAdder_138_io_co; // @[wallace.scala 67:19]
  assign FullAdder_166_io_a = FullAdder_98_io_co; // @[wallace.scala 65:18]
  assign FullAdder_166_io_b = FullAdder_99_io_co; // @[wallace.scala 66:18]
  assign FullAdder_166_io_ci = FullAdder_138_io_s; // @[wallace.scala 67:19]
  assign FullAdder_167_io_a = FullAdder_139_io_s; // @[wallace.scala 65:18]
  assign FullAdder_167_io_b = FullAdder_140_io_co; // @[wallace.scala 66:18]
  assign FullAdder_167_io_ci = FullAdder_141_io_co; // @[wallace.scala 67:19]
  assign FullAdder_168_io_a = FullAdder_102_io_co; // @[wallace.scala 65:18]
  assign FullAdder_168_io_b = FullAdder_140_io_s; // @[wallace.scala 66:18]
  assign FullAdder_168_io_ci = FullAdder_141_io_s; // @[wallace.scala 67:19]
  assign FullAdder_169_io_a = FullAdder_104_io_co; // @[wallace.scala 65:18]
  assign FullAdder_169_io_b = FullAdder_105_io_co; // @[wallace.scala 66:18]
  assign FullAdder_169_io_ci = FullAdder_142_io_s; // @[wallace.scala 67:19]
  assign FullAdder_170_io_a = FullAdder_143_io_s; // @[wallace.scala 65:18]
  assign FullAdder_170_io_b = FullAdder_144_io_co; // @[wallace.scala 66:18]
  assign FullAdder_170_io_ci = FullAdder_145_io_co; // @[wallace.scala 67:19]
  assign FullAdder_171_io_a = FullAdder_144_io_s; // @[wallace.scala 65:18]
  assign FullAdder_171_io_b = FullAdder_145_io_s; // @[wallace.scala 66:18]
  assign FullAdder_171_io_ci = FullAdder_146_io_co; // @[wallace.scala 67:19]
  assign FullAdder_172_io_a = FullAdder_111_io_co; // @[wallace.scala 65:18]
  assign FullAdder_172_io_b = FullAdder_146_io_s; // @[wallace.scala 66:18]
  assign FullAdder_172_io_ci = FullAdder_147_io_s; // @[wallace.scala 67:19]
  assign FullAdder_173_io_a = FullAdder_112_io_co; // @[wallace.scala 65:18]
  assign FullAdder_173_io_b = FullAdder_113_io_co; // @[wallace.scala 66:18]
  assign FullAdder_173_io_ci = FullAdder_148_io_s; // @[wallace.scala 67:19]
  assign FullAdder_174_io_a = FullAdder_114_io_co; // @[wallace.scala 65:18]
  assign FullAdder_174_io_b = FullAdder_115_io_co; // @[wallace.scala 66:18]
  assign FullAdder_174_io_ci = FullAdder_149_io_s; // @[wallace.scala 67:19]
  assign HalfAdder_1_io_a = FullAdder_150_io_co; // @[wallace.scala 56:18]
  assign HalfAdder_1_io_b = FullAdder_151_io_co; // @[wallace.scala 57:18]
  assign FullAdder_175_io_a = FullAdder_150_io_s; // @[wallace.scala 65:18]
  assign FullAdder_175_io_b = FullAdder_151_io_s; // @[wallace.scala 66:18]
  assign FullAdder_175_io_ci = FullAdder_152_io_co; // @[wallace.scala 67:19]
  assign FullAdder_176_io_a = FullAdder_118_io_co; // @[wallace.scala 65:18]
  assign FullAdder_176_io_b = FullAdder_152_io_s; // @[wallace.scala 66:18]
  assign FullAdder_176_io_ci = FullAdder_153_io_co; // @[wallace.scala 67:19]
  assign FullAdder_177_io_a = FullAdder_153_io_s; // @[wallace.scala 65:18]
  assign FullAdder_177_io_b = HalfAdder_io_s; // @[wallace.scala 66:18]
  assign FullAdder_177_io_ci = FullAdder_154_io_co; // @[wallace.scala 67:19]
  assign FullAdder_178_io_a = FullAdder_122_io_s; // @[wallace.scala 65:18]
  assign FullAdder_178_io_b = FullAdder_123_io_co; // @[wallace.scala 66:18]
  assign FullAdder_178_io_ci = FullAdder_156_io_co; // @[wallace.scala 67:19]
  assign FullAdder_179_io_a = FullAdder_127_io_s; // @[wallace.scala 65:18]
  assign FullAdder_179_io_b = FullAdder_128_io_co; // @[wallace.scala 66:18]
  assign FullAdder_179_io_ci = FullAdder_159_io_co; // @[wallace.scala 67:19]
  assign FullAdder_180_io_a = FullAdder_129_io_co; // @[wallace.scala 65:18]
  assign FullAdder_180_io_b = FullAdder_159_io_s; // @[wallace.scala 66:18]
  assign FullAdder_180_io_ci = FullAdder_160_io_co; // @[wallace.scala 67:19]
  assign FullAdder_181_io_a = FullAdder_130_io_co; // @[wallace.scala 65:18]
  assign FullAdder_181_io_b = FullAdder_160_io_s; // @[wallace.scala 66:18]
  assign FullAdder_181_io_ci = FullAdder_161_io_co; // @[wallace.scala 67:19]
  assign FullAdder_182_io_a = FullAdder_132_io_co; // @[wallace.scala 65:18]
  assign FullAdder_182_io_b = FullAdder_161_io_s; // @[wallace.scala 66:18]
  assign FullAdder_182_io_ci = FullAdder_162_io_co; // @[wallace.scala 67:19]
  assign FullAdder_183_io_a = FullAdder_134_io_co; // @[wallace.scala 65:18]
  assign FullAdder_183_io_b = FullAdder_135_io_co; // @[wallace.scala 66:18]
  assign FullAdder_183_io_ci = FullAdder_163_io_s; // @[wallace.scala 67:19]
  assign FullAdder_184_io_a = FullAdder_136_io_co; // @[wallace.scala 65:18]
  assign FullAdder_184_io_b = FullAdder_137_io_co; // @[wallace.scala 66:18]
  assign FullAdder_184_io_ci = FullAdder_164_io_s; // @[wallace.scala 67:19]
  assign FullAdder_185_io_a = FullAdder_139_io_co; // @[wallace.scala 65:18]
  assign FullAdder_185_io_b = FullAdder_165_io_s; // @[wallace.scala 66:18]
  assign FullAdder_185_io_ci = FullAdder_166_io_co; // @[wallace.scala 67:19]
  assign FullAdder_186_io_a = FullAdder_166_io_s; // @[wallace.scala 65:18]
  assign FullAdder_186_io_b = FullAdder_167_io_s; // @[wallace.scala 66:18]
  assign FullAdder_186_io_ci = FullAdder_168_io_co; // @[wallace.scala 67:19]
  assign FullAdder_187_io_a = FullAdder_142_io_co; // @[wallace.scala 65:18]
  assign FullAdder_187_io_b = FullAdder_143_io_co; // @[wallace.scala 66:18]
  assign FullAdder_187_io_ci = FullAdder_168_io_s; // @[wallace.scala 67:19]
  assign HalfAdder_2_io_a = FullAdder_169_io_co; // @[wallace.scala 56:18]
  assign HalfAdder_2_io_b = FullAdder_170_io_co; // @[wallace.scala 57:18]
  assign FullAdder_188_io_a = FullAdder_169_io_s; // @[wallace.scala 65:18]
  assign FullAdder_188_io_b = FullAdder_170_io_s; // @[wallace.scala 66:18]
  assign FullAdder_188_io_ci = FullAdder_171_io_co; // @[wallace.scala 67:19]
  assign FullAdder_189_io_a = FullAdder_147_io_co; // @[wallace.scala 65:18]
  assign FullAdder_189_io_b = FullAdder_171_io_s; // @[wallace.scala 66:18]
  assign FullAdder_189_io_ci = FullAdder_172_io_co; // @[wallace.scala 67:19]
  assign FullAdder_190_io_a = FullAdder_148_io_co; // @[wallace.scala 65:18]
  assign FullAdder_190_io_b = FullAdder_172_io_s; // @[wallace.scala 66:18]
  assign FullAdder_190_io_ci = FullAdder_173_io_co; // @[wallace.scala 67:19]
  assign FullAdder_191_io_a = FullAdder_149_io_co; // @[wallace.scala 65:18]
  assign FullAdder_191_io_b = FullAdder_173_io_s; // @[wallace.scala 66:18]
  assign FullAdder_191_io_ci = FullAdder_174_io_co; // @[wallace.scala 67:19]
  assign FullAdder_192_io_a = FullAdder_174_io_s; // @[wallace.scala 65:18]
  assign FullAdder_192_io_b = HalfAdder_1_io_s; // @[wallace.scala 66:18]
  assign FullAdder_192_io_ci = FullAdder_175_io_co; // @[wallace.scala 67:19]
  assign FullAdder_193_io_a = HalfAdder_io_co; // @[wallace.scala 65:18]
  assign FullAdder_193_io_b = FullAdder_176_io_s; // @[wallace.scala 66:18]
  assign FullAdder_193_io_ci = FullAdder_177_io_co; // @[wallace.scala 67:19]
  assign FullAdder_194_io_a = FullAdder_122_io_co; // @[wallace.scala 65:18]
  assign FullAdder_194_io_b = FullAdder_155_io_s; // @[wallace.scala 66:18]
  assign FullAdder_194_io_ci = FullAdder_178_io_co; // @[wallace.scala 67:19]
  assign FullAdder_195_io_a = FullAdder_162_io_s; // @[wallace.scala 65:18]
  assign FullAdder_195_io_b = FullAdder_163_io_co; // @[wallace.scala 66:18]
  assign FullAdder_195_io_ci = FullAdder_183_io_co; // @[wallace.scala 67:19]
  assign FullAdder_196_io_a = FullAdder_164_io_co; // @[wallace.scala 65:18]
  assign FullAdder_196_io_b = FullAdder_183_io_s; // @[wallace.scala 66:18]
  assign FullAdder_196_io_ci = FullAdder_184_io_co; // @[wallace.scala 67:19]
  assign FullAdder_197_io_a = FullAdder_165_io_co; // @[wallace.scala 65:18]
  assign FullAdder_197_io_b = FullAdder_184_io_s; // @[wallace.scala 66:18]
  assign FullAdder_197_io_ci = FullAdder_185_io_co; // @[wallace.scala 67:19]
  assign FullAdder_198_io_a = FullAdder_167_io_co; // @[wallace.scala 65:18]
  assign FullAdder_198_io_b = FullAdder_185_io_s; // @[wallace.scala 66:18]
  assign FullAdder_198_io_ci = FullAdder_186_io_co; // @[wallace.scala 67:19]
  assign FullAdder_199_io_a = FullAdder_186_io_s; // @[wallace.scala 65:18]
  assign FullAdder_199_io_b = FullAdder_187_io_co; // @[wallace.scala 66:18]
  assign FullAdder_199_io_ci = HalfAdder_2_io_co; // @[wallace.scala 67:19]
  assign FullAdder_200_io_a = FullAdder_187_io_s; // @[wallace.scala 65:18]
  assign FullAdder_200_io_b = HalfAdder_2_io_s; // @[wallace.scala 66:18]
  assign FullAdder_200_io_ci = FullAdder_188_io_co; // @[wallace.scala 67:19]
  assign HalfAdder_3_io_a = FullAdder_188_io_s; // @[wallace.scala 56:18]
  assign HalfAdder_3_io_b = FullAdder_189_io_co; // @[wallace.scala 57:18]
  assign HalfAdder_4_io_a = FullAdder_189_io_s; // @[wallace.scala 56:18]
  assign HalfAdder_4_io_b = FullAdder_190_io_co; // @[wallace.scala 57:18]
  assign HalfAdder_5_io_a = FullAdder_190_io_s; // @[wallace.scala 56:18]
  assign HalfAdder_5_io_b = FullAdder_191_io_co; // @[wallace.scala 57:18]
  assign FullAdder_201_io_a = HalfAdder_1_io_co; // @[wallace.scala 65:18]
  assign FullAdder_201_io_b = FullAdder_191_io_s; // @[wallace.scala 66:18]
  assign FullAdder_201_io_ci = FullAdder_192_io_co; // @[wallace.scala 67:19]
  assign FullAdder_202_io_a = FullAdder_175_io_s; // @[wallace.scala 65:18]
  assign FullAdder_202_io_b = FullAdder_176_io_co; // @[wallace.scala 66:18]
  assign FullAdder_202_io_ci = FullAdder_193_io_co; // @[wallace.scala 67:19]
  assign FullAdder_203_io_a = FullAdder_154_io_s; // @[wallace.scala 65:18]
  assign FullAdder_203_io_b = FullAdder_155_io_co; // @[wallace.scala 66:18]
  assign FullAdder_203_io_ci = FullAdder_194_io_co; // @[wallace.scala 67:19]
endmodule
module Black(
  input   io_i_pj,
  input   io_i_gj,
  input   io_i_pk,
  input   io_i_gk,
  output  io_o_g,
  output  io_o_p
);
  wire  _T = io_i_gj & io_i_pk; // @[pg.scala 26:32]
  assign io_o_g = io_i_gk | _T; // @[pg.scala 26:10]
  assign io_o_p = io_i_pk & io_i_pj; // @[pg.scala 27:10]
endmodule
module PPAdder(
  input         clock,
  input         reset,
  input  [30:0] io_augend,
  input  [30:0] io_addend,
  output [30:0] io_outs
);
  wire  PG_io_a; // @[ppadder.scala 35:20]
  wire  PG_io_b; // @[ppadder.scala 35:20]
  wire  PG_io_s; // @[ppadder.scala 35:20]
  wire  PG_io_co; // @[ppadder.scala 35:20]
  wire  PG_1_io_a; // @[ppadder.scala 35:20]
  wire  PG_1_io_b; // @[ppadder.scala 35:20]
  wire  PG_1_io_s; // @[ppadder.scala 35:20]
  wire  PG_1_io_co; // @[ppadder.scala 35:20]
  wire  PG_2_io_a; // @[ppadder.scala 35:20]
  wire  PG_2_io_b; // @[ppadder.scala 35:20]
  wire  PG_2_io_s; // @[ppadder.scala 35:20]
  wire  PG_2_io_co; // @[ppadder.scala 35:20]
  wire  PG_3_io_a; // @[ppadder.scala 35:20]
  wire  PG_3_io_b; // @[ppadder.scala 35:20]
  wire  PG_3_io_s; // @[ppadder.scala 35:20]
  wire  PG_3_io_co; // @[ppadder.scala 35:20]
  wire  PG_4_io_a; // @[ppadder.scala 35:20]
  wire  PG_4_io_b; // @[ppadder.scala 35:20]
  wire  PG_4_io_s; // @[ppadder.scala 35:20]
  wire  PG_4_io_co; // @[ppadder.scala 35:20]
  wire  PG_5_io_a; // @[ppadder.scala 35:20]
  wire  PG_5_io_b; // @[ppadder.scala 35:20]
  wire  PG_5_io_s; // @[ppadder.scala 35:20]
  wire  PG_5_io_co; // @[ppadder.scala 35:20]
  wire  PG_6_io_a; // @[ppadder.scala 35:20]
  wire  PG_6_io_b; // @[ppadder.scala 35:20]
  wire  PG_6_io_s; // @[ppadder.scala 35:20]
  wire  PG_6_io_co; // @[ppadder.scala 35:20]
  wire  PG_7_io_a; // @[ppadder.scala 35:20]
  wire  PG_7_io_b; // @[ppadder.scala 35:20]
  wire  PG_7_io_s; // @[ppadder.scala 35:20]
  wire  PG_7_io_co; // @[ppadder.scala 35:20]
  wire  PG_8_io_a; // @[ppadder.scala 35:20]
  wire  PG_8_io_b; // @[ppadder.scala 35:20]
  wire  PG_8_io_s; // @[ppadder.scala 35:20]
  wire  PG_8_io_co; // @[ppadder.scala 35:20]
  wire  PG_9_io_a; // @[ppadder.scala 35:20]
  wire  PG_9_io_b; // @[ppadder.scala 35:20]
  wire  PG_9_io_s; // @[ppadder.scala 35:20]
  wire  PG_9_io_co; // @[ppadder.scala 35:20]
  wire  PG_10_io_a; // @[ppadder.scala 35:20]
  wire  PG_10_io_b; // @[ppadder.scala 35:20]
  wire  PG_10_io_s; // @[ppadder.scala 35:20]
  wire  PG_10_io_co; // @[ppadder.scala 35:20]
  wire  PG_11_io_a; // @[ppadder.scala 35:20]
  wire  PG_11_io_b; // @[ppadder.scala 35:20]
  wire  PG_11_io_s; // @[ppadder.scala 35:20]
  wire  PG_11_io_co; // @[ppadder.scala 35:20]
  wire  PG_12_io_a; // @[ppadder.scala 35:20]
  wire  PG_12_io_b; // @[ppadder.scala 35:20]
  wire  PG_12_io_s; // @[ppadder.scala 35:20]
  wire  PG_12_io_co; // @[ppadder.scala 35:20]
  wire  PG_13_io_a; // @[ppadder.scala 35:20]
  wire  PG_13_io_b; // @[ppadder.scala 35:20]
  wire  PG_13_io_s; // @[ppadder.scala 35:20]
  wire  PG_13_io_co; // @[ppadder.scala 35:20]
  wire  PG_14_io_a; // @[ppadder.scala 35:20]
  wire  PG_14_io_b; // @[ppadder.scala 35:20]
  wire  PG_14_io_s; // @[ppadder.scala 35:20]
  wire  PG_14_io_co; // @[ppadder.scala 35:20]
  wire  PG_15_io_a; // @[ppadder.scala 35:20]
  wire  PG_15_io_b; // @[ppadder.scala 35:20]
  wire  PG_15_io_s; // @[ppadder.scala 35:20]
  wire  PG_15_io_co; // @[ppadder.scala 35:20]
  wire  PG_16_io_a; // @[ppadder.scala 35:20]
  wire  PG_16_io_b; // @[ppadder.scala 35:20]
  wire  PG_16_io_s; // @[ppadder.scala 35:20]
  wire  PG_16_io_co; // @[ppadder.scala 35:20]
  wire  PG_17_io_a; // @[ppadder.scala 35:20]
  wire  PG_17_io_b; // @[ppadder.scala 35:20]
  wire  PG_17_io_s; // @[ppadder.scala 35:20]
  wire  PG_17_io_co; // @[ppadder.scala 35:20]
  wire  PG_18_io_a; // @[ppadder.scala 35:20]
  wire  PG_18_io_b; // @[ppadder.scala 35:20]
  wire  PG_18_io_s; // @[ppadder.scala 35:20]
  wire  PG_18_io_co; // @[ppadder.scala 35:20]
  wire  PG_19_io_a; // @[ppadder.scala 35:20]
  wire  PG_19_io_b; // @[ppadder.scala 35:20]
  wire  PG_19_io_s; // @[ppadder.scala 35:20]
  wire  PG_19_io_co; // @[ppadder.scala 35:20]
  wire  PG_20_io_a; // @[ppadder.scala 35:20]
  wire  PG_20_io_b; // @[ppadder.scala 35:20]
  wire  PG_20_io_s; // @[ppadder.scala 35:20]
  wire  PG_20_io_co; // @[ppadder.scala 35:20]
  wire  PG_21_io_a; // @[ppadder.scala 35:20]
  wire  PG_21_io_b; // @[ppadder.scala 35:20]
  wire  PG_21_io_s; // @[ppadder.scala 35:20]
  wire  PG_21_io_co; // @[ppadder.scala 35:20]
  wire  PG_22_io_a; // @[ppadder.scala 35:20]
  wire  PG_22_io_b; // @[ppadder.scala 35:20]
  wire  PG_22_io_s; // @[ppadder.scala 35:20]
  wire  PG_22_io_co; // @[ppadder.scala 35:20]
  wire  PG_23_io_a; // @[ppadder.scala 35:20]
  wire  PG_23_io_b; // @[ppadder.scala 35:20]
  wire  PG_23_io_s; // @[ppadder.scala 35:20]
  wire  PG_23_io_co; // @[ppadder.scala 35:20]
  wire  PG_24_io_a; // @[ppadder.scala 35:20]
  wire  PG_24_io_b; // @[ppadder.scala 35:20]
  wire  PG_24_io_s; // @[ppadder.scala 35:20]
  wire  PG_24_io_co; // @[ppadder.scala 35:20]
  wire  PG_25_io_a; // @[ppadder.scala 35:20]
  wire  PG_25_io_b; // @[ppadder.scala 35:20]
  wire  PG_25_io_s; // @[ppadder.scala 35:20]
  wire  PG_25_io_co; // @[ppadder.scala 35:20]
  wire  PG_26_io_a; // @[ppadder.scala 35:20]
  wire  PG_26_io_b; // @[ppadder.scala 35:20]
  wire  PG_26_io_s; // @[ppadder.scala 35:20]
  wire  PG_26_io_co; // @[ppadder.scala 35:20]
  wire  PG_27_io_a; // @[ppadder.scala 35:20]
  wire  PG_27_io_b; // @[ppadder.scala 35:20]
  wire  PG_27_io_s; // @[ppadder.scala 35:20]
  wire  PG_27_io_co; // @[ppadder.scala 35:20]
  wire  PG_28_io_a; // @[ppadder.scala 35:20]
  wire  PG_28_io_b; // @[ppadder.scala 35:20]
  wire  PG_28_io_s; // @[ppadder.scala 35:20]
  wire  PG_28_io_co; // @[ppadder.scala 35:20]
  wire  PG_29_io_a; // @[ppadder.scala 35:20]
  wire  PG_29_io_b; // @[ppadder.scala 35:20]
  wire  PG_29_io_s; // @[ppadder.scala 35:20]
  wire  PG_29_io_co; // @[ppadder.scala 35:20]
  wire  PG_30_io_a; // @[ppadder.scala 35:20]
  wire  PG_30_io_b; // @[ppadder.scala 35:20]
  wire  PG_30_io_s; // @[ppadder.scala 35:20]
  wire  PG_30_io_co; // @[ppadder.scala 35:20]
  wire  Black_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_1_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_1_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_1_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_2_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_2_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_2_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_3_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_3_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_3_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_4_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_4_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_4_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_5_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_5_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_5_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_6_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_6_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_6_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_7_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_7_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_7_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_8_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_8_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_8_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_9_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_9_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_9_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_10_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_10_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_10_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_11_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_11_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_11_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_12_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_12_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_12_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_13_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_13_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_13_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_14_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_14_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_14_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_15_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_15_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_15_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_16_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_16_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_16_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_17_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_17_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_17_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_18_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_18_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_18_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_19_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_19_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_19_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_20_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_20_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_20_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_21_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_21_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_21_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_22_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_22_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_22_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_23_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_23_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_23_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_24_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_24_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_24_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_25_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_25_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_25_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_26_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_26_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_26_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_27_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_27_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_27_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_28_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_28_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_28_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_29_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_29_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_29_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_30_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_30_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_30_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_31_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_31_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_31_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_32_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_32_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_32_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_33_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_33_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_33_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_34_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_34_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_34_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_35_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_35_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_35_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_36_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_36_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_36_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_37_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_37_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_37_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_38_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_38_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_38_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_39_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_39_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_39_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_40_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_40_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_40_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_41_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_41_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_41_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_42_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_42_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_42_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_43_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_43_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_43_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_44_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_44_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_44_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_45_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_45_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_45_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_46_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_46_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_46_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_47_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_47_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_47_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_48_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_48_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_48_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_49_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_49_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_49_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_50_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_50_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_50_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_51_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_51_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_51_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_52_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_52_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_52_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_53_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_53_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_53_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_54_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_54_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_54_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_55_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_55_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_55_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_56_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_56_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_56_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_57_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_57_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_57_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_58_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_58_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_58_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_59_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_59_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_59_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_60_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_60_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_60_io_o_p; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_pj; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_gj; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_pk; // @[ppadder.scala 62:23]
  wire  Black_61_io_i_gk; // @[ppadder.scala 62:23]
  wire  Black_61_io_o_g; // @[ppadder.scala 62:23]
  wire  Black_61_io_o_p; // @[ppadder.scala 62:23]
  wire  res_0 = PG_io_s; // @[ppadder.scala 76:40]
  wire  _T_64 = ~reset; // @[ppadder.scala 77:9]
  wire  res_1 = PG_1_io_s ^ PG_io_co; // @[ppadder.scala 80:43]
  wire  res_2 = PG_2_io_s ^ Black_32_io_o_g; // @[ppadder.scala 80:43]
  wire  res_3 = PG_3_io_s ^ Black_61_io_o_g; // @[ppadder.scala 80:43]
  wire  res_4 = PG_4_io_s ^ Black_33_io_o_g; // @[ppadder.scala 80:43]
  wire  res_5 = PG_5_io_s ^ Black_59_io_o_g; // @[ppadder.scala 80:43]
  wire  res_6 = PG_6_io_s ^ Black_60_io_o_g; // @[ppadder.scala 80:43]
  wire  res_7 = PG_7_io_s ^ Black_34_io_o_g; // @[ppadder.scala 80:43]
  wire  res_8 = PG_8_io_s ^ Black_58_io_o_g; // @[ppadder.scala 80:43]
  wire  res_9 = PG_9_io_s ^ Black_57_io_o_g; // @[ppadder.scala 80:43]
  wire  res_10 = PG_10_io_s ^ Black_55_io_o_g; // @[ppadder.scala 80:43]
  wire  res_11 = PG_11_io_s ^ Black_56_io_o_g; // @[ppadder.scala 80:43]
  wire  res_12 = PG_12_io_s ^ Black_35_io_o_g; // @[ppadder.scala 80:43]
  wire  res_13 = PG_13_io_s ^ Black_54_io_o_g; // @[ppadder.scala 80:43]
  wire  res_14 = PG_14_io_s ^ Black_53_io_o_g; // @[ppadder.scala 80:43]
  wire  res_15 = PG_15_io_s ^ Black_52_io_o_g; // @[ppadder.scala 80:43]
  wire  res_16 = PG_16_io_s ^ Black_51_io_o_g; // @[ppadder.scala 80:43]
  wire  res_17 = PG_17_io_s ^ Black_36_io_o_g; // @[ppadder.scala 80:43]
  wire  res_18 = PG_18_io_s ^ Black_50_io_o_g; // @[ppadder.scala 80:43]
  wire  res_19 = PG_19_io_s ^ Black_49_io_o_g; // @[ppadder.scala 80:43]
  wire  res_20 = PG_20_io_s ^ Black_48_io_o_g; // @[ppadder.scala 80:43]
  wire  res_21 = PG_21_io_s ^ Black_47_io_o_g; // @[ppadder.scala 80:43]
  wire  res_22 = PG_22_io_s ^ Black_46_io_o_g; // @[ppadder.scala 80:43]
  wire  res_23 = PG_23_io_s ^ Black_45_io_o_g; // @[ppadder.scala 80:43]
  wire  res_24 = PG_24_io_s ^ Black_44_io_o_g; // @[ppadder.scala 80:43]
  wire  res_25 = PG_25_io_s ^ Black_43_io_o_g; // @[ppadder.scala 80:43]
  wire  res_26 = PG_26_io_s ^ Black_42_io_o_g; // @[ppadder.scala 80:43]
  wire  res_27 = PG_27_io_s ^ Black_41_io_o_g; // @[ppadder.scala 80:43]
  wire  res_28 = PG_28_io_s ^ Black_40_io_o_g; // @[ppadder.scala 80:43]
  wire  res_29 = PG_29_io_s ^ Black_39_io_o_g; // @[ppadder.scala 80:43]
  wire  res_30 = PG_30_io_s ^ Black_38_io_o_g; // @[ppadder.scala 80:43]
  wire [9:0] _T_103 = {res_30,res_29,res_28,res_27,res_26,res_25,res_24,res_23,res_22,res_21}; // @[Cat.scala 29:58]
  wire [18:0] _T_112 = {_T_103,res_20,res_19,res_18,res_17,res_16,res_15,res_14,res_13,res_12}; // @[Cat.scala 29:58]
  wire [27:0] _T_121 = {_T_112,res_11,res_10,res_9,res_8,res_7,res_6,res_5,res_4,res_3}; // @[Cat.scala 29:58]
  wire [29:0] _T_123 = {_T_121,res_2,res_1}; // @[Cat.scala 29:58]
  HalfAdder PG ( // @[ppadder.scala 35:20]
    .io_a(PG_io_a),
    .io_b(PG_io_b),
    .io_s(PG_io_s),
    .io_co(PG_io_co)
  );
  HalfAdder PG_1 ( // @[ppadder.scala 35:20]
    .io_a(PG_1_io_a),
    .io_b(PG_1_io_b),
    .io_s(PG_1_io_s),
    .io_co(PG_1_io_co)
  );
  HalfAdder PG_2 ( // @[ppadder.scala 35:20]
    .io_a(PG_2_io_a),
    .io_b(PG_2_io_b),
    .io_s(PG_2_io_s),
    .io_co(PG_2_io_co)
  );
  HalfAdder PG_3 ( // @[ppadder.scala 35:20]
    .io_a(PG_3_io_a),
    .io_b(PG_3_io_b),
    .io_s(PG_3_io_s),
    .io_co(PG_3_io_co)
  );
  HalfAdder PG_4 ( // @[ppadder.scala 35:20]
    .io_a(PG_4_io_a),
    .io_b(PG_4_io_b),
    .io_s(PG_4_io_s),
    .io_co(PG_4_io_co)
  );
  HalfAdder PG_5 ( // @[ppadder.scala 35:20]
    .io_a(PG_5_io_a),
    .io_b(PG_5_io_b),
    .io_s(PG_5_io_s),
    .io_co(PG_5_io_co)
  );
  HalfAdder PG_6 ( // @[ppadder.scala 35:20]
    .io_a(PG_6_io_a),
    .io_b(PG_6_io_b),
    .io_s(PG_6_io_s),
    .io_co(PG_6_io_co)
  );
  HalfAdder PG_7 ( // @[ppadder.scala 35:20]
    .io_a(PG_7_io_a),
    .io_b(PG_7_io_b),
    .io_s(PG_7_io_s),
    .io_co(PG_7_io_co)
  );
  HalfAdder PG_8 ( // @[ppadder.scala 35:20]
    .io_a(PG_8_io_a),
    .io_b(PG_8_io_b),
    .io_s(PG_8_io_s),
    .io_co(PG_8_io_co)
  );
  HalfAdder PG_9 ( // @[ppadder.scala 35:20]
    .io_a(PG_9_io_a),
    .io_b(PG_9_io_b),
    .io_s(PG_9_io_s),
    .io_co(PG_9_io_co)
  );
  HalfAdder PG_10 ( // @[ppadder.scala 35:20]
    .io_a(PG_10_io_a),
    .io_b(PG_10_io_b),
    .io_s(PG_10_io_s),
    .io_co(PG_10_io_co)
  );
  HalfAdder PG_11 ( // @[ppadder.scala 35:20]
    .io_a(PG_11_io_a),
    .io_b(PG_11_io_b),
    .io_s(PG_11_io_s),
    .io_co(PG_11_io_co)
  );
  HalfAdder PG_12 ( // @[ppadder.scala 35:20]
    .io_a(PG_12_io_a),
    .io_b(PG_12_io_b),
    .io_s(PG_12_io_s),
    .io_co(PG_12_io_co)
  );
  HalfAdder PG_13 ( // @[ppadder.scala 35:20]
    .io_a(PG_13_io_a),
    .io_b(PG_13_io_b),
    .io_s(PG_13_io_s),
    .io_co(PG_13_io_co)
  );
  HalfAdder PG_14 ( // @[ppadder.scala 35:20]
    .io_a(PG_14_io_a),
    .io_b(PG_14_io_b),
    .io_s(PG_14_io_s),
    .io_co(PG_14_io_co)
  );
  HalfAdder PG_15 ( // @[ppadder.scala 35:20]
    .io_a(PG_15_io_a),
    .io_b(PG_15_io_b),
    .io_s(PG_15_io_s),
    .io_co(PG_15_io_co)
  );
  HalfAdder PG_16 ( // @[ppadder.scala 35:20]
    .io_a(PG_16_io_a),
    .io_b(PG_16_io_b),
    .io_s(PG_16_io_s),
    .io_co(PG_16_io_co)
  );
  HalfAdder PG_17 ( // @[ppadder.scala 35:20]
    .io_a(PG_17_io_a),
    .io_b(PG_17_io_b),
    .io_s(PG_17_io_s),
    .io_co(PG_17_io_co)
  );
  HalfAdder PG_18 ( // @[ppadder.scala 35:20]
    .io_a(PG_18_io_a),
    .io_b(PG_18_io_b),
    .io_s(PG_18_io_s),
    .io_co(PG_18_io_co)
  );
  HalfAdder PG_19 ( // @[ppadder.scala 35:20]
    .io_a(PG_19_io_a),
    .io_b(PG_19_io_b),
    .io_s(PG_19_io_s),
    .io_co(PG_19_io_co)
  );
  HalfAdder PG_20 ( // @[ppadder.scala 35:20]
    .io_a(PG_20_io_a),
    .io_b(PG_20_io_b),
    .io_s(PG_20_io_s),
    .io_co(PG_20_io_co)
  );
  HalfAdder PG_21 ( // @[ppadder.scala 35:20]
    .io_a(PG_21_io_a),
    .io_b(PG_21_io_b),
    .io_s(PG_21_io_s),
    .io_co(PG_21_io_co)
  );
  HalfAdder PG_22 ( // @[ppadder.scala 35:20]
    .io_a(PG_22_io_a),
    .io_b(PG_22_io_b),
    .io_s(PG_22_io_s),
    .io_co(PG_22_io_co)
  );
  HalfAdder PG_23 ( // @[ppadder.scala 35:20]
    .io_a(PG_23_io_a),
    .io_b(PG_23_io_b),
    .io_s(PG_23_io_s),
    .io_co(PG_23_io_co)
  );
  HalfAdder PG_24 ( // @[ppadder.scala 35:20]
    .io_a(PG_24_io_a),
    .io_b(PG_24_io_b),
    .io_s(PG_24_io_s),
    .io_co(PG_24_io_co)
  );
  HalfAdder PG_25 ( // @[ppadder.scala 35:20]
    .io_a(PG_25_io_a),
    .io_b(PG_25_io_b),
    .io_s(PG_25_io_s),
    .io_co(PG_25_io_co)
  );
  HalfAdder PG_26 ( // @[ppadder.scala 35:20]
    .io_a(PG_26_io_a),
    .io_b(PG_26_io_b),
    .io_s(PG_26_io_s),
    .io_co(PG_26_io_co)
  );
  HalfAdder PG_27 ( // @[ppadder.scala 35:20]
    .io_a(PG_27_io_a),
    .io_b(PG_27_io_b),
    .io_s(PG_27_io_s),
    .io_co(PG_27_io_co)
  );
  HalfAdder PG_28 ( // @[ppadder.scala 35:20]
    .io_a(PG_28_io_a),
    .io_b(PG_28_io_b),
    .io_s(PG_28_io_s),
    .io_co(PG_28_io_co)
  );
  HalfAdder PG_29 ( // @[ppadder.scala 35:20]
    .io_a(PG_29_io_a),
    .io_b(PG_29_io_b),
    .io_s(PG_29_io_s),
    .io_co(PG_29_io_co)
  );
  HalfAdder PG_30 ( // @[ppadder.scala 35:20]
    .io_a(PG_30_io_a),
    .io_b(PG_30_io_b),
    .io_s(PG_30_io_s),
    .io_co(PG_30_io_co)
  );
  Black Black ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_io_i_pj),
    .io_i_gj(Black_io_i_gj),
    .io_i_pk(Black_io_i_pk),
    .io_i_gk(Black_io_i_gk),
    .io_o_g(Black_io_o_g),
    .io_o_p(Black_io_o_p)
  );
  Black Black_1 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_1_io_i_pj),
    .io_i_gj(Black_1_io_i_gj),
    .io_i_pk(Black_1_io_i_pk),
    .io_i_gk(Black_1_io_i_gk),
    .io_o_g(Black_1_io_o_g),
    .io_o_p(Black_1_io_o_p)
  );
  Black Black_2 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_2_io_i_pj),
    .io_i_gj(Black_2_io_i_gj),
    .io_i_pk(Black_2_io_i_pk),
    .io_i_gk(Black_2_io_i_gk),
    .io_o_g(Black_2_io_o_g),
    .io_o_p(Black_2_io_o_p)
  );
  Black Black_3 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_3_io_i_pj),
    .io_i_gj(Black_3_io_i_gj),
    .io_i_pk(Black_3_io_i_pk),
    .io_i_gk(Black_3_io_i_gk),
    .io_o_g(Black_3_io_o_g),
    .io_o_p(Black_3_io_o_p)
  );
  Black Black_4 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_4_io_i_pj),
    .io_i_gj(Black_4_io_i_gj),
    .io_i_pk(Black_4_io_i_pk),
    .io_i_gk(Black_4_io_i_gk),
    .io_o_g(Black_4_io_o_g),
    .io_o_p(Black_4_io_o_p)
  );
  Black Black_5 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_5_io_i_pj),
    .io_i_gj(Black_5_io_i_gj),
    .io_i_pk(Black_5_io_i_pk),
    .io_i_gk(Black_5_io_i_gk),
    .io_o_g(Black_5_io_o_g),
    .io_o_p(Black_5_io_o_p)
  );
  Black Black_6 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_6_io_i_pj),
    .io_i_gj(Black_6_io_i_gj),
    .io_i_pk(Black_6_io_i_pk),
    .io_i_gk(Black_6_io_i_gk),
    .io_o_g(Black_6_io_o_g),
    .io_o_p(Black_6_io_o_p)
  );
  Black Black_7 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_7_io_i_pj),
    .io_i_gj(Black_7_io_i_gj),
    .io_i_pk(Black_7_io_i_pk),
    .io_i_gk(Black_7_io_i_gk),
    .io_o_g(Black_7_io_o_g),
    .io_o_p(Black_7_io_o_p)
  );
  Black Black_8 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_8_io_i_pj),
    .io_i_gj(Black_8_io_i_gj),
    .io_i_pk(Black_8_io_i_pk),
    .io_i_gk(Black_8_io_i_gk),
    .io_o_g(Black_8_io_o_g),
    .io_o_p(Black_8_io_o_p)
  );
  Black Black_9 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_9_io_i_pj),
    .io_i_gj(Black_9_io_i_gj),
    .io_i_pk(Black_9_io_i_pk),
    .io_i_gk(Black_9_io_i_gk),
    .io_o_g(Black_9_io_o_g),
    .io_o_p(Black_9_io_o_p)
  );
  Black Black_10 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_10_io_i_pj),
    .io_i_gj(Black_10_io_i_gj),
    .io_i_pk(Black_10_io_i_pk),
    .io_i_gk(Black_10_io_i_gk),
    .io_o_g(Black_10_io_o_g),
    .io_o_p(Black_10_io_o_p)
  );
  Black Black_11 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_11_io_i_pj),
    .io_i_gj(Black_11_io_i_gj),
    .io_i_pk(Black_11_io_i_pk),
    .io_i_gk(Black_11_io_i_gk),
    .io_o_g(Black_11_io_o_g),
    .io_o_p(Black_11_io_o_p)
  );
  Black Black_12 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_12_io_i_pj),
    .io_i_gj(Black_12_io_i_gj),
    .io_i_pk(Black_12_io_i_pk),
    .io_i_gk(Black_12_io_i_gk),
    .io_o_g(Black_12_io_o_g),
    .io_o_p(Black_12_io_o_p)
  );
  Black Black_13 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_13_io_i_pj),
    .io_i_gj(Black_13_io_i_gj),
    .io_i_pk(Black_13_io_i_pk),
    .io_i_gk(Black_13_io_i_gk),
    .io_o_g(Black_13_io_o_g),
    .io_o_p(Black_13_io_o_p)
  );
  Black Black_14 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_14_io_i_pj),
    .io_i_gj(Black_14_io_i_gj),
    .io_i_pk(Black_14_io_i_pk),
    .io_i_gk(Black_14_io_i_gk),
    .io_o_g(Black_14_io_o_g),
    .io_o_p(Black_14_io_o_p)
  );
  Black Black_15 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_15_io_i_pj),
    .io_i_gj(Black_15_io_i_gj),
    .io_i_pk(Black_15_io_i_pk),
    .io_i_gk(Black_15_io_i_gk),
    .io_o_g(Black_15_io_o_g),
    .io_o_p(Black_15_io_o_p)
  );
  Black Black_16 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_16_io_i_pj),
    .io_i_gj(Black_16_io_i_gj),
    .io_i_pk(Black_16_io_i_pk),
    .io_i_gk(Black_16_io_i_gk),
    .io_o_g(Black_16_io_o_g),
    .io_o_p(Black_16_io_o_p)
  );
  Black Black_17 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_17_io_i_pj),
    .io_i_gj(Black_17_io_i_gj),
    .io_i_pk(Black_17_io_i_pk),
    .io_i_gk(Black_17_io_i_gk),
    .io_o_g(Black_17_io_o_g),
    .io_o_p(Black_17_io_o_p)
  );
  Black Black_18 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_18_io_i_pj),
    .io_i_gj(Black_18_io_i_gj),
    .io_i_pk(Black_18_io_i_pk),
    .io_i_gk(Black_18_io_i_gk),
    .io_o_g(Black_18_io_o_g),
    .io_o_p(Black_18_io_o_p)
  );
  Black Black_19 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_19_io_i_pj),
    .io_i_gj(Black_19_io_i_gj),
    .io_i_pk(Black_19_io_i_pk),
    .io_i_gk(Black_19_io_i_gk),
    .io_o_g(Black_19_io_o_g),
    .io_o_p(Black_19_io_o_p)
  );
  Black Black_20 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_20_io_i_pj),
    .io_i_gj(Black_20_io_i_gj),
    .io_i_pk(Black_20_io_i_pk),
    .io_i_gk(Black_20_io_i_gk),
    .io_o_g(Black_20_io_o_g),
    .io_o_p(Black_20_io_o_p)
  );
  Black Black_21 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_21_io_i_pj),
    .io_i_gj(Black_21_io_i_gj),
    .io_i_pk(Black_21_io_i_pk),
    .io_i_gk(Black_21_io_i_gk),
    .io_o_g(Black_21_io_o_g),
    .io_o_p(Black_21_io_o_p)
  );
  Black Black_22 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_22_io_i_pj),
    .io_i_gj(Black_22_io_i_gj),
    .io_i_pk(Black_22_io_i_pk),
    .io_i_gk(Black_22_io_i_gk),
    .io_o_g(Black_22_io_o_g),
    .io_o_p(Black_22_io_o_p)
  );
  Black Black_23 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_23_io_i_pj),
    .io_i_gj(Black_23_io_i_gj),
    .io_i_pk(Black_23_io_i_pk),
    .io_i_gk(Black_23_io_i_gk),
    .io_o_g(Black_23_io_o_g),
    .io_o_p(Black_23_io_o_p)
  );
  Black Black_24 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_24_io_i_pj),
    .io_i_gj(Black_24_io_i_gj),
    .io_i_pk(Black_24_io_i_pk),
    .io_i_gk(Black_24_io_i_gk),
    .io_o_g(Black_24_io_o_g),
    .io_o_p(Black_24_io_o_p)
  );
  Black Black_25 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_25_io_i_pj),
    .io_i_gj(Black_25_io_i_gj),
    .io_i_pk(Black_25_io_i_pk),
    .io_i_gk(Black_25_io_i_gk),
    .io_o_g(Black_25_io_o_g),
    .io_o_p(Black_25_io_o_p)
  );
  Black Black_26 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_26_io_i_pj),
    .io_i_gj(Black_26_io_i_gj),
    .io_i_pk(Black_26_io_i_pk),
    .io_i_gk(Black_26_io_i_gk),
    .io_o_g(Black_26_io_o_g),
    .io_o_p(Black_26_io_o_p)
  );
  Black Black_27 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_27_io_i_pj),
    .io_i_gj(Black_27_io_i_gj),
    .io_i_pk(Black_27_io_i_pk),
    .io_i_gk(Black_27_io_i_gk),
    .io_o_g(Black_27_io_o_g),
    .io_o_p(Black_27_io_o_p)
  );
  Black Black_28 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_28_io_i_pj),
    .io_i_gj(Black_28_io_i_gj),
    .io_i_pk(Black_28_io_i_pk),
    .io_i_gk(Black_28_io_i_gk),
    .io_o_g(Black_28_io_o_g),
    .io_o_p(Black_28_io_o_p)
  );
  Black Black_29 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_29_io_i_pj),
    .io_i_gj(Black_29_io_i_gj),
    .io_i_pk(Black_29_io_i_pk),
    .io_i_gk(Black_29_io_i_gk),
    .io_o_g(Black_29_io_o_g),
    .io_o_p(Black_29_io_o_p)
  );
  Black Black_30 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_30_io_i_pj),
    .io_i_gj(Black_30_io_i_gj),
    .io_i_pk(Black_30_io_i_pk),
    .io_i_gk(Black_30_io_i_gk),
    .io_o_g(Black_30_io_o_g),
    .io_o_p(Black_30_io_o_p)
  );
  Black Black_31 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_31_io_i_pj),
    .io_i_gj(Black_31_io_i_gj),
    .io_i_pk(Black_31_io_i_pk),
    .io_i_gk(Black_31_io_i_gk),
    .io_o_g(Black_31_io_o_g),
    .io_o_p(Black_31_io_o_p)
  );
  Black Black_32 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_32_io_i_pj),
    .io_i_gj(Black_32_io_i_gj),
    .io_i_pk(Black_32_io_i_pk),
    .io_i_gk(Black_32_io_i_gk),
    .io_o_g(Black_32_io_o_g),
    .io_o_p(Black_32_io_o_p)
  );
  Black Black_33 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_33_io_i_pj),
    .io_i_gj(Black_33_io_i_gj),
    .io_i_pk(Black_33_io_i_pk),
    .io_i_gk(Black_33_io_i_gk),
    .io_o_g(Black_33_io_o_g),
    .io_o_p(Black_33_io_o_p)
  );
  Black Black_34 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_34_io_i_pj),
    .io_i_gj(Black_34_io_i_gj),
    .io_i_pk(Black_34_io_i_pk),
    .io_i_gk(Black_34_io_i_gk),
    .io_o_g(Black_34_io_o_g),
    .io_o_p(Black_34_io_o_p)
  );
  Black Black_35 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_35_io_i_pj),
    .io_i_gj(Black_35_io_i_gj),
    .io_i_pk(Black_35_io_i_pk),
    .io_i_gk(Black_35_io_i_gk),
    .io_o_g(Black_35_io_o_g),
    .io_o_p(Black_35_io_o_p)
  );
  Black Black_36 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_36_io_i_pj),
    .io_i_gj(Black_36_io_i_gj),
    .io_i_pk(Black_36_io_i_pk),
    .io_i_gk(Black_36_io_i_gk),
    .io_o_g(Black_36_io_o_g),
    .io_o_p(Black_36_io_o_p)
  );
  Black Black_37 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_37_io_i_pj),
    .io_i_gj(Black_37_io_i_gj),
    .io_i_pk(Black_37_io_i_pk),
    .io_i_gk(Black_37_io_i_gk),
    .io_o_g(Black_37_io_o_g),
    .io_o_p(Black_37_io_o_p)
  );
  Black Black_38 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_38_io_i_pj),
    .io_i_gj(Black_38_io_i_gj),
    .io_i_pk(Black_38_io_i_pk),
    .io_i_gk(Black_38_io_i_gk),
    .io_o_g(Black_38_io_o_g),
    .io_o_p(Black_38_io_o_p)
  );
  Black Black_39 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_39_io_i_pj),
    .io_i_gj(Black_39_io_i_gj),
    .io_i_pk(Black_39_io_i_pk),
    .io_i_gk(Black_39_io_i_gk),
    .io_o_g(Black_39_io_o_g),
    .io_o_p(Black_39_io_o_p)
  );
  Black Black_40 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_40_io_i_pj),
    .io_i_gj(Black_40_io_i_gj),
    .io_i_pk(Black_40_io_i_pk),
    .io_i_gk(Black_40_io_i_gk),
    .io_o_g(Black_40_io_o_g),
    .io_o_p(Black_40_io_o_p)
  );
  Black Black_41 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_41_io_i_pj),
    .io_i_gj(Black_41_io_i_gj),
    .io_i_pk(Black_41_io_i_pk),
    .io_i_gk(Black_41_io_i_gk),
    .io_o_g(Black_41_io_o_g),
    .io_o_p(Black_41_io_o_p)
  );
  Black Black_42 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_42_io_i_pj),
    .io_i_gj(Black_42_io_i_gj),
    .io_i_pk(Black_42_io_i_pk),
    .io_i_gk(Black_42_io_i_gk),
    .io_o_g(Black_42_io_o_g),
    .io_o_p(Black_42_io_o_p)
  );
  Black Black_43 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_43_io_i_pj),
    .io_i_gj(Black_43_io_i_gj),
    .io_i_pk(Black_43_io_i_pk),
    .io_i_gk(Black_43_io_i_gk),
    .io_o_g(Black_43_io_o_g),
    .io_o_p(Black_43_io_o_p)
  );
  Black Black_44 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_44_io_i_pj),
    .io_i_gj(Black_44_io_i_gj),
    .io_i_pk(Black_44_io_i_pk),
    .io_i_gk(Black_44_io_i_gk),
    .io_o_g(Black_44_io_o_g),
    .io_o_p(Black_44_io_o_p)
  );
  Black Black_45 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_45_io_i_pj),
    .io_i_gj(Black_45_io_i_gj),
    .io_i_pk(Black_45_io_i_pk),
    .io_i_gk(Black_45_io_i_gk),
    .io_o_g(Black_45_io_o_g),
    .io_o_p(Black_45_io_o_p)
  );
  Black Black_46 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_46_io_i_pj),
    .io_i_gj(Black_46_io_i_gj),
    .io_i_pk(Black_46_io_i_pk),
    .io_i_gk(Black_46_io_i_gk),
    .io_o_g(Black_46_io_o_g),
    .io_o_p(Black_46_io_o_p)
  );
  Black Black_47 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_47_io_i_pj),
    .io_i_gj(Black_47_io_i_gj),
    .io_i_pk(Black_47_io_i_pk),
    .io_i_gk(Black_47_io_i_gk),
    .io_o_g(Black_47_io_o_g),
    .io_o_p(Black_47_io_o_p)
  );
  Black Black_48 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_48_io_i_pj),
    .io_i_gj(Black_48_io_i_gj),
    .io_i_pk(Black_48_io_i_pk),
    .io_i_gk(Black_48_io_i_gk),
    .io_o_g(Black_48_io_o_g),
    .io_o_p(Black_48_io_o_p)
  );
  Black Black_49 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_49_io_i_pj),
    .io_i_gj(Black_49_io_i_gj),
    .io_i_pk(Black_49_io_i_pk),
    .io_i_gk(Black_49_io_i_gk),
    .io_o_g(Black_49_io_o_g),
    .io_o_p(Black_49_io_o_p)
  );
  Black Black_50 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_50_io_i_pj),
    .io_i_gj(Black_50_io_i_gj),
    .io_i_pk(Black_50_io_i_pk),
    .io_i_gk(Black_50_io_i_gk),
    .io_o_g(Black_50_io_o_g),
    .io_o_p(Black_50_io_o_p)
  );
  Black Black_51 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_51_io_i_pj),
    .io_i_gj(Black_51_io_i_gj),
    .io_i_pk(Black_51_io_i_pk),
    .io_i_gk(Black_51_io_i_gk),
    .io_o_g(Black_51_io_o_g),
    .io_o_p(Black_51_io_o_p)
  );
  Black Black_52 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_52_io_i_pj),
    .io_i_gj(Black_52_io_i_gj),
    .io_i_pk(Black_52_io_i_pk),
    .io_i_gk(Black_52_io_i_gk),
    .io_o_g(Black_52_io_o_g),
    .io_o_p(Black_52_io_o_p)
  );
  Black Black_53 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_53_io_i_pj),
    .io_i_gj(Black_53_io_i_gj),
    .io_i_pk(Black_53_io_i_pk),
    .io_i_gk(Black_53_io_i_gk),
    .io_o_g(Black_53_io_o_g),
    .io_o_p(Black_53_io_o_p)
  );
  Black Black_54 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_54_io_i_pj),
    .io_i_gj(Black_54_io_i_gj),
    .io_i_pk(Black_54_io_i_pk),
    .io_i_gk(Black_54_io_i_gk),
    .io_o_g(Black_54_io_o_g),
    .io_o_p(Black_54_io_o_p)
  );
  Black Black_55 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_55_io_i_pj),
    .io_i_gj(Black_55_io_i_gj),
    .io_i_pk(Black_55_io_i_pk),
    .io_i_gk(Black_55_io_i_gk),
    .io_o_g(Black_55_io_o_g),
    .io_o_p(Black_55_io_o_p)
  );
  Black Black_56 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_56_io_i_pj),
    .io_i_gj(Black_56_io_i_gj),
    .io_i_pk(Black_56_io_i_pk),
    .io_i_gk(Black_56_io_i_gk),
    .io_o_g(Black_56_io_o_g),
    .io_o_p(Black_56_io_o_p)
  );
  Black Black_57 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_57_io_i_pj),
    .io_i_gj(Black_57_io_i_gj),
    .io_i_pk(Black_57_io_i_pk),
    .io_i_gk(Black_57_io_i_gk),
    .io_o_g(Black_57_io_o_g),
    .io_o_p(Black_57_io_o_p)
  );
  Black Black_58 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_58_io_i_pj),
    .io_i_gj(Black_58_io_i_gj),
    .io_i_pk(Black_58_io_i_pk),
    .io_i_gk(Black_58_io_i_gk),
    .io_o_g(Black_58_io_o_g),
    .io_o_p(Black_58_io_o_p)
  );
  Black Black_59 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_59_io_i_pj),
    .io_i_gj(Black_59_io_i_gj),
    .io_i_pk(Black_59_io_i_pk),
    .io_i_gk(Black_59_io_i_gk),
    .io_o_g(Black_59_io_o_g),
    .io_o_p(Black_59_io_o_p)
  );
  Black Black_60 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_60_io_i_pj),
    .io_i_gj(Black_60_io_i_gj),
    .io_i_pk(Black_60_io_i_pk),
    .io_i_gk(Black_60_io_i_gk),
    .io_o_g(Black_60_io_o_g),
    .io_o_p(Black_60_io_o_p)
  );
  Black Black_61 ( // @[ppadder.scala 62:23]
    .io_i_pj(Black_61_io_i_pj),
    .io_i_gj(Black_61_io_i_gj),
    .io_i_pk(Black_61_io_i_pk),
    .io_i_gk(Black_61_io_i_gk),
    .io_o_g(Black_61_io_o_g),
    .io_o_p(Black_61_io_o_p)
  );
  assign io_outs = {_T_123,res_0}; // @[ppadder.scala 84:11]
  assign PG_io_a = io_augend[0]; // @[ppadder.scala 36:15]
  assign PG_io_b = io_addend[0]; // @[ppadder.scala 37:15]
  assign PG_1_io_a = io_augend[1]; // @[ppadder.scala 36:15]
  assign PG_1_io_b = io_addend[1]; // @[ppadder.scala 37:15]
  assign PG_2_io_a = io_augend[2]; // @[ppadder.scala 36:15]
  assign PG_2_io_b = io_addend[2]; // @[ppadder.scala 37:15]
  assign PG_3_io_a = io_augend[3]; // @[ppadder.scala 36:15]
  assign PG_3_io_b = io_addend[3]; // @[ppadder.scala 37:15]
  assign PG_4_io_a = io_augend[4]; // @[ppadder.scala 36:15]
  assign PG_4_io_b = io_addend[4]; // @[ppadder.scala 37:15]
  assign PG_5_io_a = io_augend[5]; // @[ppadder.scala 36:15]
  assign PG_5_io_b = io_addend[5]; // @[ppadder.scala 37:15]
  assign PG_6_io_a = io_augend[6]; // @[ppadder.scala 36:15]
  assign PG_6_io_b = io_addend[6]; // @[ppadder.scala 37:15]
  assign PG_7_io_a = io_augend[7]; // @[ppadder.scala 36:15]
  assign PG_7_io_b = io_addend[7]; // @[ppadder.scala 37:15]
  assign PG_8_io_a = io_augend[8]; // @[ppadder.scala 36:15]
  assign PG_8_io_b = io_addend[8]; // @[ppadder.scala 37:15]
  assign PG_9_io_a = io_augend[9]; // @[ppadder.scala 36:15]
  assign PG_9_io_b = io_addend[9]; // @[ppadder.scala 37:15]
  assign PG_10_io_a = io_augend[10]; // @[ppadder.scala 36:15]
  assign PG_10_io_b = io_addend[10]; // @[ppadder.scala 37:15]
  assign PG_11_io_a = io_augend[11]; // @[ppadder.scala 36:15]
  assign PG_11_io_b = io_addend[11]; // @[ppadder.scala 37:15]
  assign PG_12_io_a = io_augend[12]; // @[ppadder.scala 36:15]
  assign PG_12_io_b = io_addend[12]; // @[ppadder.scala 37:15]
  assign PG_13_io_a = io_augend[13]; // @[ppadder.scala 36:15]
  assign PG_13_io_b = io_addend[13]; // @[ppadder.scala 37:15]
  assign PG_14_io_a = io_augend[14]; // @[ppadder.scala 36:15]
  assign PG_14_io_b = io_addend[14]; // @[ppadder.scala 37:15]
  assign PG_15_io_a = io_augend[15]; // @[ppadder.scala 36:15]
  assign PG_15_io_b = io_addend[15]; // @[ppadder.scala 37:15]
  assign PG_16_io_a = io_augend[16]; // @[ppadder.scala 36:15]
  assign PG_16_io_b = io_addend[16]; // @[ppadder.scala 37:15]
  assign PG_17_io_a = io_augend[17]; // @[ppadder.scala 36:15]
  assign PG_17_io_b = io_addend[17]; // @[ppadder.scala 37:15]
  assign PG_18_io_a = io_augend[18]; // @[ppadder.scala 36:15]
  assign PG_18_io_b = io_addend[18]; // @[ppadder.scala 37:15]
  assign PG_19_io_a = io_augend[19]; // @[ppadder.scala 36:15]
  assign PG_19_io_b = io_addend[19]; // @[ppadder.scala 37:15]
  assign PG_20_io_a = io_augend[20]; // @[ppadder.scala 36:15]
  assign PG_20_io_b = io_addend[20]; // @[ppadder.scala 37:15]
  assign PG_21_io_a = io_augend[21]; // @[ppadder.scala 36:15]
  assign PG_21_io_b = io_addend[21]; // @[ppadder.scala 37:15]
  assign PG_22_io_a = io_augend[22]; // @[ppadder.scala 36:15]
  assign PG_22_io_b = io_addend[22]; // @[ppadder.scala 37:15]
  assign PG_23_io_a = io_augend[23]; // @[ppadder.scala 36:15]
  assign PG_23_io_b = io_addend[23]; // @[ppadder.scala 37:15]
  assign PG_24_io_a = io_augend[24]; // @[ppadder.scala 36:15]
  assign PG_24_io_b = io_addend[24]; // @[ppadder.scala 37:15]
  assign PG_25_io_a = io_augend[25]; // @[ppadder.scala 36:15]
  assign PG_25_io_b = io_addend[25]; // @[ppadder.scala 37:15]
  assign PG_26_io_a = io_augend[26]; // @[ppadder.scala 36:15]
  assign PG_26_io_b = io_addend[26]; // @[ppadder.scala 37:15]
  assign PG_27_io_a = io_augend[27]; // @[ppadder.scala 36:15]
  assign PG_27_io_b = io_addend[27]; // @[ppadder.scala 37:15]
  assign PG_28_io_a = io_augend[28]; // @[ppadder.scala 36:15]
  assign PG_28_io_b = io_addend[28]; // @[ppadder.scala 37:15]
  assign PG_29_io_a = io_augend[29]; // @[ppadder.scala 36:15]
  assign PG_29_io_b = io_addend[29]; // @[ppadder.scala 37:15]
  assign PG_30_io_a = io_augend[30]; // @[ppadder.scala 36:15]
  assign PG_30_io_b = io_addend[30]; // @[ppadder.scala 37:15]
  assign Black_io_i_pj = PG_26_io_s; // @[ppadder.scala 66:19]
  assign Black_io_i_gj = PG_26_io_co; // @[ppadder.scala 65:19]
  assign Black_io_i_pk = PG_27_io_s; // @[ppadder.scala 64:19]
  assign Black_io_i_gk = PG_27_io_co; // @[ppadder.scala 63:19]
  assign Black_1_io_i_pj = Black_io_o_p; // @[ppadder.scala 66:19]
  assign Black_1_io_i_gj = Black_io_o_g; // @[ppadder.scala 65:19]
  assign Black_1_io_i_pk = PG_28_io_s; // @[ppadder.scala 64:19]
  assign Black_1_io_i_gk = PG_28_io_co; // @[ppadder.scala 63:19]
  assign Black_2_io_i_pj = Black_1_io_o_p; // @[ppadder.scala 66:19]
  assign Black_2_io_i_gj = Black_1_io_o_g; // @[ppadder.scala 65:19]
  assign Black_2_io_i_pk = PG_29_io_s; // @[ppadder.scala 64:19]
  assign Black_2_io_i_gk = PG_29_io_co; // @[ppadder.scala 63:19]
  assign Black_3_io_i_pj = Black_2_io_o_p; // @[ppadder.scala 66:19]
  assign Black_3_io_i_gj = Black_2_io_o_g; // @[ppadder.scala 65:19]
  assign Black_3_io_i_pk = PG_30_io_s; // @[ppadder.scala 64:19]
  assign Black_3_io_i_gk = PG_30_io_co; // @[ppadder.scala 63:19]
  assign Black_4_io_i_pj = PG_22_io_s; // @[ppadder.scala 66:19]
  assign Black_4_io_i_gj = PG_22_io_co; // @[ppadder.scala 65:19]
  assign Black_4_io_i_pk = PG_23_io_s; // @[ppadder.scala 64:19]
  assign Black_4_io_i_gk = PG_23_io_co; // @[ppadder.scala 63:19]
  assign Black_5_io_i_pj = Black_4_io_o_p; // @[ppadder.scala 66:19]
  assign Black_5_io_i_gj = Black_4_io_o_g; // @[ppadder.scala 65:19]
  assign Black_5_io_i_pk = PG_24_io_s; // @[ppadder.scala 64:19]
  assign Black_5_io_i_gk = PG_24_io_co; // @[ppadder.scala 63:19]
  assign Black_6_io_i_pj = Black_5_io_o_p; // @[ppadder.scala 66:19]
  assign Black_6_io_i_gj = Black_5_io_o_g; // @[ppadder.scala 65:19]
  assign Black_6_io_i_pk = PG_25_io_s; // @[ppadder.scala 64:19]
  assign Black_6_io_i_gk = PG_25_io_co; // @[ppadder.scala 63:19]
  assign Black_7_io_i_pj = PG_20_io_s; // @[ppadder.scala 66:19]
  assign Black_7_io_i_gj = PG_20_io_co; // @[ppadder.scala 65:19]
  assign Black_7_io_i_pk = PG_21_io_s; // @[ppadder.scala 64:19]
  assign Black_7_io_i_gk = PG_21_io_co; // @[ppadder.scala 63:19]
  assign Black_8_io_i_pj = PG_17_io_s; // @[ppadder.scala 66:19]
  assign Black_8_io_i_gj = PG_17_io_co; // @[ppadder.scala 65:19]
  assign Black_8_io_i_pk = PG_18_io_s; // @[ppadder.scala 64:19]
  assign Black_8_io_i_gk = PG_18_io_co; // @[ppadder.scala 63:19]
  assign Black_9_io_i_pj = Black_8_io_o_p; // @[ppadder.scala 66:19]
  assign Black_9_io_i_gj = Black_8_io_o_g; // @[ppadder.scala 65:19]
  assign Black_9_io_i_pk = PG_19_io_s; // @[ppadder.scala 64:19]
  assign Black_9_io_i_gk = PG_19_io_co; // @[ppadder.scala 63:19]
  assign Black_10_io_i_pj = Black_9_io_o_p; // @[ppadder.scala 66:19]
  assign Black_10_io_i_gj = Black_9_io_o_g; // @[ppadder.scala 65:19]
  assign Black_10_io_i_pk = Black_7_io_o_p; // @[ppadder.scala 64:19]
  assign Black_10_io_i_gk = Black_7_io_o_g; // @[ppadder.scala 63:19]
  assign Black_11_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_11_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_11_io_i_pk = Black_6_io_o_p; // @[ppadder.scala 64:19]
  assign Black_11_io_i_gk = Black_6_io_o_g; // @[ppadder.scala 63:19]
  assign Black_12_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_12_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_12_io_i_pk = Black_3_io_o_p; // @[ppadder.scala 64:19]
  assign Black_12_io_i_gk = Black_3_io_o_g; // @[ppadder.scala 63:19]
  assign Black_13_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_13_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_13_io_i_pk = Black_2_io_o_p; // @[ppadder.scala 64:19]
  assign Black_13_io_i_gk = Black_2_io_o_g; // @[ppadder.scala 63:19]
  assign Black_14_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_14_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_14_io_i_pk = Black_1_io_o_p; // @[ppadder.scala 64:19]
  assign Black_14_io_i_gk = Black_1_io_o_g; // @[ppadder.scala 63:19]
  assign Black_15_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_15_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_15_io_i_pk = Black_io_o_p; // @[ppadder.scala 64:19]
  assign Black_15_io_i_gk = Black_io_o_g; // @[ppadder.scala 63:19]
  assign Black_16_io_i_pj = Black_11_io_o_p; // @[ppadder.scala 66:19]
  assign Black_16_io_i_gj = Black_11_io_o_g; // @[ppadder.scala 65:19]
  assign Black_16_io_i_pk = PG_26_io_s; // @[ppadder.scala 64:19]
  assign Black_16_io_i_gk = PG_26_io_co; // @[ppadder.scala 63:19]
  assign Black_17_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_17_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_17_io_i_pk = Black_5_io_o_p; // @[ppadder.scala 64:19]
  assign Black_17_io_i_gk = Black_5_io_o_g; // @[ppadder.scala 63:19]
  assign Black_18_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_18_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_18_io_i_pk = Black_4_io_o_p; // @[ppadder.scala 64:19]
  assign Black_18_io_i_gk = Black_4_io_o_g; // @[ppadder.scala 63:19]
  assign Black_19_io_i_pj = Black_10_io_o_p; // @[ppadder.scala 66:19]
  assign Black_19_io_i_gj = Black_10_io_o_g; // @[ppadder.scala 65:19]
  assign Black_19_io_i_pk = PG_22_io_s; // @[ppadder.scala 64:19]
  assign Black_19_io_i_gk = PG_22_io_co; // @[ppadder.scala 63:19]
  assign Black_20_io_i_pj = Black_9_io_o_p; // @[ppadder.scala 66:19]
  assign Black_20_io_i_gj = Black_9_io_o_g; // @[ppadder.scala 65:19]
  assign Black_20_io_i_pk = PG_20_io_s; // @[ppadder.scala 64:19]
  assign Black_20_io_i_gk = PG_20_io_co; // @[ppadder.scala 63:19]
  assign Black_21_io_i_pj = PG_12_io_s; // @[ppadder.scala 66:19]
  assign Black_21_io_i_gj = PG_12_io_co; // @[ppadder.scala 65:19]
  assign Black_21_io_i_pk = PG_13_io_s; // @[ppadder.scala 64:19]
  assign Black_21_io_i_gk = PG_13_io_co; // @[ppadder.scala 63:19]
  assign Black_22_io_i_pj = Black_21_io_o_p; // @[ppadder.scala 66:19]
  assign Black_22_io_i_gj = Black_21_io_o_g; // @[ppadder.scala 65:19]
  assign Black_22_io_i_pk = PG_14_io_s; // @[ppadder.scala 64:19]
  assign Black_22_io_i_gk = PG_14_io_co; // @[ppadder.scala 63:19]
  assign Black_23_io_i_pj = Black_22_io_o_p; // @[ppadder.scala 66:19]
  assign Black_23_io_i_gj = Black_22_io_o_g; // @[ppadder.scala 65:19]
  assign Black_23_io_i_pk = PG_15_io_s; // @[ppadder.scala 64:19]
  assign Black_23_io_i_gk = PG_15_io_co; // @[ppadder.scala 63:19]
  assign Black_24_io_i_pj = Black_23_io_o_p; // @[ppadder.scala 66:19]
  assign Black_24_io_i_gj = Black_23_io_o_g; // @[ppadder.scala 65:19]
  assign Black_24_io_i_pk = PG_16_io_s; // @[ppadder.scala 64:19]
  assign Black_24_io_i_gk = PG_16_io_co; // @[ppadder.scala 63:19]
  assign Black_25_io_i_pj = PG_10_io_s; // @[ppadder.scala 66:19]
  assign Black_25_io_i_gj = PG_10_io_co; // @[ppadder.scala 65:19]
  assign Black_25_io_i_pk = PG_11_io_s; // @[ppadder.scala 64:19]
  assign Black_25_io_i_gk = PG_11_io_co; // @[ppadder.scala 63:19]
  assign Black_26_io_i_pj = PG_7_io_s; // @[ppadder.scala 66:19]
  assign Black_26_io_i_gj = PG_7_io_co; // @[ppadder.scala 65:19]
  assign Black_26_io_i_pk = PG_8_io_s; // @[ppadder.scala 64:19]
  assign Black_26_io_i_gk = PG_8_io_co; // @[ppadder.scala 63:19]
  assign Black_27_io_i_pj = Black_26_io_o_p; // @[ppadder.scala 66:19]
  assign Black_27_io_i_gj = Black_26_io_o_g; // @[ppadder.scala 65:19]
  assign Black_27_io_i_pk = PG_9_io_s; // @[ppadder.scala 64:19]
  assign Black_27_io_i_gk = PG_9_io_co; // @[ppadder.scala 63:19]
  assign Black_28_io_i_pj = Black_27_io_o_p; // @[ppadder.scala 66:19]
  assign Black_28_io_i_gj = Black_27_io_o_g; // @[ppadder.scala 65:19]
  assign Black_28_io_i_pk = Black_25_io_o_p; // @[ppadder.scala 64:19]
  assign Black_28_io_i_gk = Black_25_io_o_g; // @[ppadder.scala 63:19]
  assign Black_29_io_i_pj = PG_5_io_s; // @[ppadder.scala 66:19]
  assign Black_29_io_i_gj = PG_5_io_co; // @[ppadder.scala 65:19]
  assign Black_29_io_i_pk = PG_6_io_s; // @[ppadder.scala 64:19]
  assign Black_29_io_i_gk = PG_6_io_co; // @[ppadder.scala 63:19]
  assign Black_30_io_i_pj = PG_4_io_s; // @[ppadder.scala 66:19]
  assign Black_30_io_i_gj = PG_4_io_co; // @[ppadder.scala 65:19]
  assign Black_30_io_i_pk = Black_29_io_o_p; // @[ppadder.scala 64:19]
  assign Black_30_io_i_gk = Black_29_io_o_g; // @[ppadder.scala 63:19]
  assign Black_31_io_i_pj = PG_2_io_s; // @[ppadder.scala 66:19]
  assign Black_31_io_i_gj = PG_2_io_co; // @[ppadder.scala 65:19]
  assign Black_31_io_i_pk = PG_3_io_s; // @[ppadder.scala 64:19]
  assign Black_31_io_i_gk = PG_3_io_co; // @[ppadder.scala 63:19]
  assign Black_32_io_i_pj = PG_io_s; // @[ppadder.scala 66:19]
  assign Black_32_io_i_gj = PG_io_co; // @[ppadder.scala 65:19]
  assign Black_32_io_i_pk = PG_1_io_s; // @[ppadder.scala 64:19]
  assign Black_32_io_i_gk = PG_1_io_co; // @[ppadder.scala 63:19]
  assign Black_33_io_i_pj = Black_32_io_o_p; // @[ppadder.scala 66:19]
  assign Black_33_io_i_gj = Black_32_io_o_g; // @[ppadder.scala 65:19]
  assign Black_33_io_i_pk = Black_31_io_o_p; // @[ppadder.scala 64:19]
  assign Black_33_io_i_gk = Black_31_io_o_g; // @[ppadder.scala 63:19]
  assign Black_34_io_i_pj = Black_33_io_o_p; // @[ppadder.scala 66:19]
  assign Black_34_io_i_gj = Black_33_io_o_g; // @[ppadder.scala 65:19]
  assign Black_34_io_i_pk = Black_30_io_o_p; // @[ppadder.scala 64:19]
  assign Black_34_io_i_gk = Black_30_io_o_g; // @[ppadder.scala 63:19]
  assign Black_35_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_35_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_35_io_i_pk = Black_28_io_o_p; // @[ppadder.scala 64:19]
  assign Black_35_io_i_gk = Black_28_io_o_g; // @[ppadder.scala 63:19]
  assign Black_36_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_36_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_36_io_i_pk = Black_24_io_o_p; // @[ppadder.scala 64:19]
  assign Black_36_io_i_gk = Black_24_io_o_g; // @[ppadder.scala 63:19]
  assign Black_37_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_37_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_37_io_i_pk = Black_12_io_o_p; // @[ppadder.scala 64:19]
  assign Black_37_io_i_gk = Black_12_io_o_g; // @[ppadder.scala 63:19]
  assign Black_38_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_38_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_38_io_i_pk = Black_13_io_o_p; // @[ppadder.scala 64:19]
  assign Black_38_io_i_gk = Black_13_io_o_g; // @[ppadder.scala 63:19]
  assign Black_39_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_39_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_39_io_i_pk = Black_14_io_o_p; // @[ppadder.scala 64:19]
  assign Black_39_io_i_gk = Black_14_io_o_g; // @[ppadder.scala 63:19]
  assign Black_40_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_40_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_40_io_i_pk = Black_15_io_o_p; // @[ppadder.scala 64:19]
  assign Black_40_io_i_gk = Black_15_io_o_g; // @[ppadder.scala 63:19]
  assign Black_41_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_41_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_41_io_i_pk = Black_16_io_o_p; // @[ppadder.scala 64:19]
  assign Black_41_io_i_gk = Black_16_io_o_g; // @[ppadder.scala 63:19]
  assign Black_42_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_42_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_42_io_i_pk = Black_11_io_o_p; // @[ppadder.scala 64:19]
  assign Black_42_io_i_gk = Black_11_io_o_g; // @[ppadder.scala 63:19]
  assign Black_43_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_43_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_43_io_i_pk = Black_17_io_o_p; // @[ppadder.scala 64:19]
  assign Black_43_io_i_gk = Black_17_io_o_g; // @[ppadder.scala 63:19]
  assign Black_44_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_44_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_44_io_i_pk = Black_18_io_o_p; // @[ppadder.scala 64:19]
  assign Black_44_io_i_gk = Black_18_io_o_g; // @[ppadder.scala 63:19]
  assign Black_45_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_45_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_45_io_i_pk = Black_19_io_o_p; // @[ppadder.scala 64:19]
  assign Black_45_io_i_gk = Black_19_io_o_g; // @[ppadder.scala 63:19]
  assign Black_46_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_46_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_46_io_i_pk = Black_10_io_o_p; // @[ppadder.scala 64:19]
  assign Black_46_io_i_gk = Black_10_io_o_g; // @[ppadder.scala 63:19]
  assign Black_47_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_47_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_47_io_i_pk = Black_20_io_o_p; // @[ppadder.scala 64:19]
  assign Black_47_io_i_gk = Black_20_io_o_g; // @[ppadder.scala 63:19]
  assign Black_48_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_48_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_48_io_i_pk = Black_9_io_o_p; // @[ppadder.scala 64:19]
  assign Black_48_io_i_gk = Black_9_io_o_g; // @[ppadder.scala 63:19]
  assign Black_49_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_49_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_49_io_i_pk = Black_8_io_o_p; // @[ppadder.scala 64:19]
  assign Black_49_io_i_gk = Black_8_io_o_g; // @[ppadder.scala 63:19]
  assign Black_50_io_i_pj = Black_36_io_o_p; // @[ppadder.scala 66:19]
  assign Black_50_io_i_gj = Black_36_io_o_g; // @[ppadder.scala 65:19]
  assign Black_50_io_i_pk = PG_17_io_s; // @[ppadder.scala 64:19]
  assign Black_50_io_i_gk = PG_17_io_co; // @[ppadder.scala 63:19]
  assign Black_51_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_51_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_51_io_i_pk = Black_23_io_o_p; // @[ppadder.scala 64:19]
  assign Black_51_io_i_gk = Black_23_io_o_g; // @[ppadder.scala 63:19]
  assign Black_52_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_52_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_52_io_i_pk = Black_22_io_o_p; // @[ppadder.scala 64:19]
  assign Black_52_io_i_gk = Black_22_io_o_g; // @[ppadder.scala 63:19]
  assign Black_53_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_53_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_53_io_i_pk = Black_21_io_o_p; // @[ppadder.scala 64:19]
  assign Black_53_io_i_gk = Black_21_io_o_g; // @[ppadder.scala 63:19]
  assign Black_54_io_i_pj = Black_35_io_o_p; // @[ppadder.scala 66:19]
  assign Black_54_io_i_gj = Black_35_io_o_g; // @[ppadder.scala 65:19]
  assign Black_54_io_i_pk = PG_12_io_s; // @[ppadder.scala 64:19]
  assign Black_54_io_i_gk = PG_12_io_co; // @[ppadder.scala 63:19]
  assign Black_55_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_55_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_55_io_i_pk = Black_27_io_o_p; // @[ppadder.scala 64:19]
  assign Black_55_io_i_gk = Black_27_io_o_g; // @[ppadder.scala 63:19]
  assign Black_56_io_i_pj = Black_55_io_o_p; // @[ppadder.scala 66:19]
  assign Black_56_io_i_gj = Black_55_io_o_g; // @[ppadder.scala 65:19]
  assign Black_56_io_i_pk = PG_10_io_s; // @[ppadder.scala 64:19]
  assign Black_56_io_i_gk = PG_10_io_co; // @[ppadder.scala 63:19]
  assign Black_57_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_57_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_57_io_i_pk = Black_26_io_o_p; // @[ppadder.scala 64:19]
  assign Black_57_io_i_gk = Black_26_io_o_g; // @[ppadder.scala 63:19]
  assign Black_58_io_i_pj = Black_34_io_o_p; // @[ppadder.scala 66:19]
  assign Black_58_io_i_gj = Black_34_io_o_g; // @[ppadder.scala 65:19]
  assign Black_58_io_i_pk = PG_7_io_s; // @[ppadder.scala 64:19]
  assign Black_58_io_i_gk = PG_7_io_co; // @[ppadder.scala 63:19]
  assign Black_59_io_i_pj = Black_33_io_o_p; // @[ppadder.scala 66:19]
  assign Black_59_io_i_gj = Black_33_io_o_g; // @[ppadder.scala 65:19]
  assign Black_59_io_i_pk = PG_4_io_s; // @[ppadder.scala 64:19]
  assign Black_59_io_i_gk = PG_4_io_co; // @[ppadder.scala 63:19]
  assign Black_60_io_i_pj = Black_59_io_o_p; // @[ppadder.scala 66:19]
  assign Black_60_io_i_gj = Black_59_io_o_g; // @[ppadder.scala 65:19]
  assign Black_60_io_i_pk = PG_5_io_s; // @[ppadder.scala 64:19]
  assign Black_60_io_i_gk = PG_5_io_co; // @[ppadder.scala 63:19]
  assign Black_61_io_i_pj = Black_32_io_o_p; // @[ppadder.scala 66:19]
  assign Black_61_io_i_gj = Black_32_io_o_g; // @[ppadder.scala 65:19]
  assign Black_61_io_i_pk = PG_2_io_s; // @[ppadder.scala 64:19]
  assign Black_61_io_i_gk = PG_2_io_co; // @[ppadder.scala 63:19]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_64) begin
          $fwrite(32'h80000002,"res(0) = %d\n",res_0); // @[ppadder.scala 77:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MAC(
  input         clock,
  input         reset,
  input  [15:0] io_multiplicand,
  input  [15:0] io_multiplier,
  input  [30:0] io_addend,
  output [30:0] io_outs
);
  wire [15:0] pp_io_multiplicand; // @[mac.scala 28:18]
  wire [15:0] pp_io_multiplier; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_0; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_1; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_2; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_3; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_4; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_5; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_6; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_7; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_8; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_9; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_10; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_11; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_12; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_13; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_14; // @[mac.scala 28:18]
  wire [15:0] pp_io_outs_15; // @[mac.scala 28:18]
  wire [15:0] wt_io_pp_0; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_1; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_2; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_3; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_4; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_5; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_6; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_7; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_8; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_9; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_10; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_11; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_12; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_13; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_14; // @[mac.scala 32:18]
  wire [15:0] wt_io_pp_15; // @[mac.scala 32:18]
  wire [31:0] wt_io_augend; // @[mac.scala 32:18]
  wire [31:0] wt_io_addend; // @[mac.scala 32:18]
  wire  ppa1_clock; // @[mac.scala 35:20]
  wire  ppa1_reset; // @[mac.scala 35:20]
  wire [30:0] ppa1_io_augend; // @[mac.scala 35:20]
  wire [30:0] ppa1_io_addend; // @[mac.scala 35:20]
  wire [30:0] ppa1_io_outs; // @[mac.scala 35:20]
  wire  ppa2_clock; // @[mac.scala 39:20]
  wire  ppa2_reset; // @[mac.scala 39:20]
  wire [30:0] ppa2_io_augend; // @[mac.scala 39:20]
  wire [30:0] ppa2_io_addend; // @[mac.scala 39:20]
  wire [30:0] ppa2_io_outs; // @[mac.scala 39:20]
  PartialProd pp ( // @[mac.scala 28:18]
    .io_multiplicand(pp_io_multiplicand),
    .io_multiplier(pp_io_multiplier),
    .io_outs_0(pp_io_outs_0),
    .io_outs_1(pp_io_outs_1),
    .io_outs_2(pp_io_outs_2),
    .io_outs_3(pp_io_outs_3),
    .io_outs_4(pp_io_outs_4),
    .io_outs_5(pp_io_outs_5),
    .io_outs_6(pp_io_outs_6),
    .io_outs_7(pp_io_outs_7),
    .io_outs_8(pp_io_outs_8),
    .io_outs_9(pp_io_outs_9),
    .io_outs_10(pp_io_outs_10),
    .io_outs_11(pp_io_outs_11),
    .io_outs_12(pp_io_outs_12),
    .io_outs_13(pp_io_outs_13),
    .io_outs_14(pp_io_outs_14),
    .io_outs_15(pp_io_outs_15)
  );
  Wallace wt ( // @[mac.scala 32:18]
    .io_pp_0(wt_io_pp_0),
    .io_pp_1(wt_io_pp_1),
    .io_pp_2(wt_io_pp_2),
    .io_pp_3(wt_io_pp_3),
    .io_pp_4(wt_io_pp_4),
    .io_pp_5(wt_io_pp_5),
    .io_pp_6(wt_io_pp_6),
    .io_pp_7(wt_io_pp_7),
    .io_pp_8(wt_io_pp_8),
    .io_pp_9(wt_io_pp_9),
    .io_pp_10(wt_io_pp_10),
    .io_pp_11(wt_io_pp_11),
    .io_pp_12(wt_io_pp_12),
    .io_pp_13(wt_io_pp_13),
    .io_pp_14(wt_io_pp_14),
    .io_pp_15(wt_io_pp_15),
    .io_augend(wt_io_augend),
    .io_addend(wt_io_addend)
  );
  PPAdder ppa1 ( // @[mac.scala 35:20]
    .clock(ppa1_clock),
    .reset(ppa1_reset),
    .io_augend(ppa1_io_augend),
    .io_addend(ppa1_io_addend),
    .io_outs(ppa1_io_outs)
  );
  PPAdder ppa2 ( // @[mac.scala 39:20]
    .clock(ppa2_clock),
    .reset(ppa2_reset),
    .io_augend(ppa2_io_augend),
    .io_addend(ppa2_io_addend),
    .io_outs(ppa2_io_outs)
  );
  assign io_outs = ppa2_io_outs; // @[mac.scala 43:11]
  assign pp_io_multiplicand = io_multiplicand; // @[mac.scala 29:22]
  assign pp_io_multiplier = io_multiplier; // @[mac.scala 30:20]
  assign wt_io_pp_0 = pp_io_outs_0; // @[mac.scala 33:12]
  assign wt_io_pp_1 = pp_io_outs_1; // @[mac.scala 33:12]
  assign wt_io_pp_2 = pp_io_outs_2; // @[mac.scala 33:12]
  assign wt_io_pp_3 = pp_io_outs_3; // @[mac.scala 33:12]
  assign wt_io_pp_4 = pp_io_outs_4; // @[mac.scala 33:12]
  assign wt_io_pp_5 = pp_io_outs_5; // @[mac.scala 33:12]
  assign wt_io_pp_6 = pp_io_outs_6; // @[mac.scala 33:12]
  assign wt_io_pp_7 = pp_io_outs_7; // @[mac.scala 33:12]
  assign wt_io_pp_8 = pp_io_outs_8; // @[mac.scala 33:12]
  assign wt_io_pp_9 = pp_io_outs_9; // @[mac.scala 33:12]
  assign wt_io_pp_10 = pp_io_outs_10; // @[mac.scala 33:12]
  assign wt_io_pp_11 = pp_io_outs_11; // @[mac.scala 33:12]
  assign wt_io_pp_12 = pp_io_outs_12; // @[mac.scala 33:12]
  assign wt_io_pp_13 = pp_io_outs_13; // @[mac.scala 33:12]
  assign wt_io_pp_14 = pp_io_outs_14; // @[mac.scala 33:12]
  assign wt_io_pp_15 = pp_io_outs_15; // @[mac.scala 33:12]
  assign ppa1_clock = clock;
  assign ppa1_reset = reset;
  assign ppa1_io_augend = wt_io_augend[30:0]; // @[mac.scala 36:18]
  assign ppa1_io_addend = wt_io_addend[30:0]; // @[mac.scala 37:18]
  assign ppa2_clock = clock;
  assign ppa2_reset = reset;
  assign ppa2_io_augend = ppa1_io_outs; // @[mac.scala 40:18]
  assign ppa2_io_addend = io_addend; // @[mac.scala 41:18]
endmodule
